magic
tech gf180mcuD
magscale 1 10
timestamp 1699643579
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 22094 38274 22146 38286
rect 19506 38222 19518 38274
rect 19570 38222 19582 38274
rect 22094 38210 22146 38222
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 21298 37998 21310 38050
rect 21362 37998 21374 38050
rect 16942 37938 16994 37950
rect 16942 37874 16994 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18510 37490 18562 37502
rect 18510 37426 18562 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 17490 37214 17502 37266
rect 17554 37214 17566 37266
rect 20850 37214 20862 37266
rect 20914 37214 20926 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 40238 36370 40290 36382
rect 40238 36306 40290 36318
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 20738 27134 20750 27186
rect 20802 27134 20814 27186
rect 21646 27074 21698 27086
rect 17938 27022 17950 27074
rect 18002 27022 18014 27074
rect 21646 27010 21698 27022
rect 18610 26910 18622 26962
rect 18674 26910 18686 26962
rect 21298 26910 21310 26962
rect 21362 26910 21374 26962
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 17390 26402 17442 26414
rect 17390 26338 17442 26350
rect 13906 26238 13918 26290
rect 13970 26238 13982 26290
rect 26562 26238 26574 26290
rect 26626 26238 26638 26290
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 17950 26178 18002 26190
rect 14690 26126 14702 26178
rect 14754 26126 14766 26178
rect 16818 26126 16830 26178
rect 16882 26126 16894 26178
rect 17950 26114 18002 26126
rect 20974 26178 21026 26190
rect 20974 26114 21026 26126
rect 24334 26178 24386 26190
rect 24334 26114 24386 26126
rect 26238 26178 26290 26190
rect 27346 26126 27358 26178
rect 27410 26126 27422 26178
rect 29474 26126 29486 26178
rect 29538 26126 29550 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 26238 26114 26290 26126
rect 17502 26066 17554 26078
rect 17502 26002 17554 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 27358 25730 27410 25742
rect 27358 25666 27410 25678
rect 1934 25618 1986 25630
rect 40014 25618 40066 25630
rect 16594 25566 16606 25618
rect 16658 25566 16670 25618
rect 22530 25566 22542 25618
rect 22594 25566 22606 25618
rect 1934 25554 1986 25566
rect 40014 25554 40066 25566
rect 27470 25506 27522 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 13458 25454 13470 25506
rect 13522 25454 13534 25506
rect 19394 25454 19406 25506
rect 19458 25454 19470 25506
rect 25330 25454 25342 25506
rect 25394 25454 25406 25506
rect 29250 25454 29262 25506
rect 29314 25454 29326 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 27470 25442 27522 25454
rect 13806 25394 13858 25406
rect 27918 25394 27970 25406
rect 18722 25342 18734 25394
rect 18786 25342 18798 25394
rect 24658 25342 24670 25394
rect 24722 25342 24734 25394
rect 13806 25330 13858 25342
rect 27918 25330 27970 25342
rect 28030 25394 28082 25406
rect 28030 25330 28082 25342
rect 13694 25282 13746 25294
rect 13694 25218 13746 25230
rect 19966 25282 20018 25294
rect 19966 25218 20018 25230
rect 25902 25282 25954 25294
rect 25902 25218 25954 25230
rect 26350 25282 26402 25294
rect 26350 25218 26402 25230
rect 27358 25282 27410 25294
rect 27358 25218 27410 25230
rect 27694 25282 27746 25294
rect 29474 25230 29486 25282
rect 29538 25230 29550 25282
rect 27694 25218 27746 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 15262 24946 15314 24958
rect 15262 24882 15314 24894
rect 15374 24946 15426 24958
rect 15374 24882 15426 24894
rect 17614 24946 17666 24958
rect 17614 24882 17666 24894
rect 17726 24946 17778 24958
rect 17726 24882 17778 24894
rect 18846 24946 18898 24958
rect 18846 24882 18898 24894
rect 19294 24946 19346 24958
rect 19294 24882 19346 24894
rect 20414 24946 20466 24958
rect 20414 24882 20466 24894
rect 24782 24946 24834 24958
rect 24782 24882 24834 24894
rect 18958 24834 19010 24846
rect 13906 24782 13918 24834
rect 13970 24782 13982 24834
rect 18958 24770 19010 24782
rect 24558 24834 24610 24846
rect 24558 24770 24610 24782
rect 15486 24722 15538 24734
rect 17502 24722 17554 24734
rect 14690 24670 14702 24722
rect 14754 24670 14766 24722
rect 15026 24670 15038 24722
rect 15090 24670 15102 24722
rect 15698 24670 15710 24722
rect 15762 24670 15774 24722
rect 15486 24658 15538 24670
rect 17502 24658 17554 24670
rect 17838 24722 17890 24734
rect 17838 24658 17890 24670
rect 17950 24722 18002 24734
rect 19742 24722 19794 24734
rect 19506 24670 19518 24722
rect 19570 24670 19582 24722
rect 17950 24658 18002 24670
rect 19742 24658 19794 24670
rect 20078 24722 20130 24734
rect 20078 24658 20130 24670
rect 20302 24722 20354 24734
rect 20974 24722 21026 24734
rect 24446 24722 24498 24734
rect 20626 24670 20638 24722
rect 20690 24670 20702 24722
rect 21186 24670 21198 24722
rect 21250 24670 21262 24722
rect 25554 24670 25566 24722
rect 25618 24670 25630 24722
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 20302 24658 20354 24670
rect 20974 24658 21026 24670
rect 24446 24658 24498 24670
rect 11778 24558 11790 24610
rect 11842 24558 11854 24610
rect 21970 24558 21982 24610
rect 22034 24558 22046 24610
rect 24098 24558 24110 24610
rect 24162 24558 24174 24610
rect 26338 24558 26350 24610
rect 26402 24558 26414 24610
rect 28466 24558 28478 24610
rect 28530 24558 28542 24610
rect 18846 24498 18898 24510
rect 18846 24434 18898 24446
rect 19630 24498 19682 24510
rect 19630 24434 19682 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 13470 24162 13522 24174
rect 13470 24098 13522 24110
rect 27022 24162 27074 24174
rect 27022 24098 27074 24110
rect 1934 24050 1986 24062
rect 1934 23986 1986 23998
rect 18622 24050 18674 24062
rect 40014 24050 40066 24062
rect 23538 23998 23550 24050
rect 23602 23998 23614 24050
rect 18622 23986 18674 23998
rect 40014 23986 40066 23998
rect 18734 23938 18786 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 13794 23886 13806 23938
rect 13858 23886 13870 23938
rect 18734 23874 18786 23886
rect 18958 23938 19010 23950
rect 27134 23938 27186 23950
rect 19170 23886 19182 23938
rect 19234 23886 19246 23938
rect 19394 23886 19406 23938
rect 19458 23886 19470 23938
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 18958 23874 19010 23886
rect 27134 23874 27186 23886
rect 28142 23938 28194 23950
rect 28142 23874 28194 23886
rect 28478 23938 28530 23950
rect 28478 23874 28530 23886
rect 29374 23938 29426 23950
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 29374 23874 29426 23886
rect 18510 23826 18562 23838
rect 18510 23762 18562 23774
rect 27022 23826 27074 23838
rect 27022 23762 27074 23774
rect 28366 23826 28418 23838
rect 28366 23762 28418 23774
rect 13582 23714 13634 23726
rect 13582 23650 13634 23662
rect 14926 23714 14978 23726
rect 14926 23650 14978 23662
rect 29038 23714 29090 23726
rect 29038 23650 29090 23662
rect 29262 23714 29314 23726
rect 29262 23650 29314 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 14926 23378 14978 23390
rect 14926 23314 14978 23326
rect 15150 23378 15202 23390
rect 15150 23314 15202 23326
rect 15934 23378 15986 23390
rect 15934 23314 15986 23326
rect 21758 23378 21810 23390
rect 21758 23314 21810 23326
rect 21870 23378 21922 23390
rect 21870 23314 21922 23326
rect 23102 23378 23154 23390
rect 23102 23314 23154 23326
rect 26798 23378 26850 23390
rect 26798 23314 26850 23326
rect 15486 23266 15538 23278
rect 21982 23266 22034 23278
rect 13682 23214 13694 23266
rect 13746 23214 13758 23266
rect 21074 23214 21086 23266
rect 21138 23214 21150 23266
rect 22754 23214 22766 23266
rect 22818 23214 22830 23266
rect 15486 23202 15538 23214
rect 21982 23202 22034 23214
rect 15038 23154 15090 23166
rect 14466 23102 14478 23154
rect 14530 23102 14542 23154
rect 15038 23090 15090 23102
rect 15262 23154 15314 23166
rect 20638 23154 20690 23166
rect 22430 23154 22482 23166
rect 20402 23102 20414 23154
rect 20466 23102 20478 23154
rect 21298 23102 21310 23154
rect 21362 23102 21374 23154
rect 23650 23102 23662 23154
rect 23714 23102 23726 23154
rect 24098 23102 24110 23154
rect 24162 23102 24174 23154
rect 27122 23102 27134 23154
rect 27186 23102 27198 23154
rect 15262 23090 15314 23102
rect 20638 23090 20690 23102
rect 22430 23090 22482 23102
rect 19742 23042 19794 23054
rect 11554 22990 11566 23042
rect 11618 22990 11630 23042
rect 19742 22978 19794 22990
rect 24222 23042 24274 23054
rect 27906 22990 27918 23042
rect 27970 22990 27982 23042
rect 30034 22990 30046 23042
rect 30098 22990 30110 23042
rect 24222 22978 24274 22990
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 15486 22594 15538 22606
rect 15486 22530 15538 22542
rect 18734 22594 18786 22606
rect 21646 22594 21698 22606
rect 21298 22542 21310 22594
rect 21362 22542 21374 22594
rect 18734 22530 18786 22542
rect 21646 22530 21698 22542
rect 22318 22594 22370 22606
rect 22318 22530 22370 22542
rect 27918 22594 27970 22606
rect 27918 22530 27970 22542
rect 1934 22482 1986 22494
rect 1934 22418 1986 22430
rect 21870 22482 21922 22494
rect 21870 22418 21922 22430
rect 24558 22482 24610 22494
rect 24558 22418 24610 22430
rect 14030 22370 14082 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 14030 22306 14082 22318
rect 14254 22370 14306 22382
rect 24334 22370 24386 22382
rect 15474 22318 15486 22370
rect 15538 22318 15550 22370
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 17826 22318 17838 22370
rect 17890 22318 17902 22370
rect 14254 22306 14306 22318
rect 24334 22306 24386 22318
rect 28030 22370 28082 22382
rect 28030 22306 28082 22318
rect 12686 22258 12738 22270
rect 12686 22194 12738 22206
rect 12910 22258 12962 22270
rect 12910 22194 12962 22206
rect 14142 22258 14194 22270
rect 14142 22194 14194 22206
rect 14590 22258 14642 22270
rect 14590 22194 14642 22206
rect 15150 22258 15202 22270
rect 15150 22194 15202 22206
rect 16942 22258 16994 22270
rect 16942 22194 16994 22206
rect 17278 22258 17330 22270
rect 17278 22194 17330 22206
rect 18062 22258 18114 22270
rect 18062 22194 18114 22206
rect 18398 22258 18450 22270
rect 18398 22194 18450 22206
rect 18846 22258 18898 22270
rect 18846 22194 18898 22206
rect 22206 22258 22258 22270
rect 23650 22206 23662 22258
rect 23714 22206 23726 22258
rect 24098 22206 24110 22258
rect 24162 22206 24174 22258
rect 22206 22194 22258 22206
rect 12798 22146 12850 22158
rect 12798 22082 12850 22094
rect 18174 22146 18226 22158
rect 18174 22082 18226 22094
rect 18622 22146 18674 22158
rect 18622 22082 18674 22094
rect 22318 22146 22370 22158
rect 22318 22082 22370 22094
rect 27918 22146 27970 22158
rect 27918 22082 27970 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 16606 21810 16658 21822
rect 16606 21746 16658 21758
rect 17726 21810 17778 21822
rect 17726 21746 17778 21758
rect 19630 21810 19682 21822
rect 19630 21746 19682 21758
rect 22766 21810 22818 21822
rect 22766 21746 22818 21758
rect 19742 21698 19794 21710
rect 13122 21646 13134 21698
rect 13186 21646 13198 21698
rect 17378 21646 17390 21698
rect 17442 21646 17454 21698
rect 19170 21646 19182 21698
rect 19234 21646 19246 21698
rect 19742 21634 19794 21646
rect 20638 21698 20690 21710
rect 22990 21698 23042 21710
rect 24670 21698 24722 21710
rect 27806 21698 27858 21710
rect 21522 21646 21534 21698
rect 21586 21646 21598 21698
rect 22194 21646 22206 21698
rect 22258 21646 22270 21698
rect 23762 21646 23774 21698
rect 23826 21646 23838 21698
rect 24210 21646 24222 21698
rect 24274 21646 24286 21698
rect 25218 21646 25230 21698
rect 25282 21646 25294 21698
rect 20638 21634 20690 21646
rect 22990 21634 23042 21646
rect 24670 21634 24722 21646
rect 27806 21634 27858 21646
rect 14366 21586 14418 21598
rect 23102 21586 23154 21598
rect 13906 21534 13918 21586
rect 13970 21534 13982 21586
rect 16818 21534 16830 21586
rect 16882 21534 16894 21586
rect 18386 21534 18398 21586
rect 18450 21534 18462 21586
rect 18722 21534 18734 21586
rect 18786 21534 18798 21586
rect 19954 21534 19966 21586
rect 20018 21534 20030 21586
rect 20178 21534 20190 21586
rect 20242 21534 20254 21586
rect 21746 21534 21758 21586
rect 21810 21534 21822 21586
rect 22418 21534 22430 21586
rect 22482 21534 22494 21586
rect 14366 21522 14418 21534
rect 23102 21522 23154 21534
rect 24446 21586 24498 21598
rect 24446 21522 24498 21534
rect 25566 21586 25618 21598
rect 25566 21522 25618 21534
rect 27582 21586 27634 21598
rect 27582 21522 27634 21534
rect 27918 21586 27970 21598
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 27918 21522 27970 21534
rect 19182 21474 19234 21486
rect 10994 21422 11006 21474
rect 11058 21422 11070 21474
rect 19182 21410 19234 21422
rect 16494 21362 16546 21374
rect 16494 21298 16546 21310
rect 20526 21362 20578 21374
rect 20526 21298 20578 21310
rect 40014 21362 40066 21374
rect 40014 21298 40066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 19406 21026 19458 21038
rect 19406 20962 19458 20974
rect 1934 20914 1986 20926
rect 16382 20914 16434 20926
rect 16034 20862 16046 20914
rect 16098 20862 16110 20914
rect 1934 20850 1986 20862
rect 16382 20850 16434 20862
rect 17950 20914 18002 20926
rect 23538 20862 23550 20914
rect 23602 20862 23614 20914
rect 17950 20850 18002 20862
rect 14926 20802 14978 20814
rect 16718 20802 16770 20814
rect 4162 20750 4174 20802
rect 4226 20750 4238 20802
rect 15250 20750 15262 20802
rect 15314 20750 15326 20802
rect 19058 20750 19070 20802
rect 19122 20750 19134 20802
rect 19954 20750 19966 20802
rect 20018 20750 20030 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 14926 20738 14978 20750
rect 16718 20738 16770 20750
rect 15486 20690 15538 20702
rect 15486 20626 15538 20638
rect 16158 20690 16210 20702
rect 16158 20626 16210 20638
rect 17166 20690 17218 20702
rect 20414 20690 20466 20702
rect 19730 20638 19742 20690
rect 19794 20638 19806 20690
rect 17166 20626 17218 20638
rect 20414 20626 20466 20638
rect 20526 20690 20578 20702
rect 20526 20626 20578 20638
rect 15598 20578 15650 20590
rect 15598 20514 15650 20526
rect 16830 20578 16882 20590
rect 16830 20514 16882 20526
rect 16942 20578 16994 20590
rect 16942 20514 16994 20526
rect 17838 20578 17890 20590
rect 17838 20514 17890 20526
rect 18062 20578 18114 20590
rect 18062 20514 18114 20526
rect 18286 20578 18338 20590
rect 18286 20514 18338 20526
rect 19294 20578 19346 20590
rect 19294 20514 19346 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14590 20242 14642 20254
rect 18958 20242 19010 20254
rect 18610 20190 18622 20242
rect 18674 20190 18686 20242
rect 22418 20190 22430 20242
rect 22482 20190 22494 20242
rect 23090 20190 23102 20242
rect 23154 20190 23166 20242
rect 14590 20178 14642 20190
rect 18958 20178 19010 20190
rect 15486 20130 15538 20142
rect 15486 20066 15538 20078
rect 16046 20130 16098 20142
rect 16046 20066 16098 20078
rect 19406 20130 19458 20142
rect 19406 20066 19458 20078
rect 19630 20130 19682 20142
rect 19630 20066 19682 20078
rect 19966 20130 20018 20142
rect 19966 20066 20018 20078
rect 21086 20130 21138 20142
rect 21086 20066 21138 20078
rect 21982 20130 22034 20142
rect 25342 20130 25394 20142
rect 29598 20130 29650 20142
rect 24434 20078 24446 20130
rect 24498 20078 24510 20130
rect 28914 20078 28926 20130
rect 28978 20078 28990 20130
rect 21982 20066 22034 20078
rect 25342 20066 25394 20078
rect 29598 20066 29650 20078
rect 29710 20130 29762 20142
rect 29710 20066 29762 20078
rect 14814 20018 14866 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 14242 19966 14254 20018
rect 14306 19966 14318 20018
rect 14814 19954 14866 19966
rect 15262 20018 15314 20030
rect 15262 19954 15314 19966
rect 15710 20018 15762 20030
rect 15710 19954 15762 19966
rect 19294 20018 19346 20030
rect 19294 19954 19346 19966
rect 19854 20018 19906 20030
rect 19854 19954 19906 19966
rect 21422 20018 21474 20030
rect 21422 19954 21474 19966
rect 21534 20018 21586 20030
rect 21534 19954 21586 19966
rect 21870 20018 21922 20030
rect 21870 19954 21922 19966
rect 22206 20018 22258 20030
rect 22206 19954 22258 19966
rect 22766 20018 22818 20030
rect 23314 19966 23326 20018
rect 23378 19966 23390 20018
rect 24210 19966 24222 20018
rect 24274 19966 24286 20018
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 29138 19966 29150 20018
rect 29202 19966 29214 20018
rect 22766 19954 22818 19966
rect 14702 19906 14754 19918
rect 11330 19854 11342 19906
rect 11394 19854 11406 19906
rect 13458 19854 13470 19906
rect 13522 19854 13534 19906
rect 14702 19842 14754 19854
rect 15598 19906 15650 19918
rect 26450 19854 26462 19906
rect 26514 19854 26526 19906
rect 28578 19854 28590 19906
rect 28642 19854 28654 19906
rect 15598 19842 15650 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 19966 19794 20018 19806
rect 19966 19730 20018 19742
rect 29710 19794 29762 19806
rect 29710 19730 29762 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 13694 19458 13746 19470
rect 13694 19394 13746 19406
rect 14030 19458 14082 19470
rect 15038 19458 15090 19470
rect 14242 19406 14254 19458
rect 14306 19455 14318 19458
rect 14690 19455 14702 19458
rect 14306 19409 14702 19455
rect 14306 19406 14318 19409
rect 14690 19406 14702 19409
rect 14754 19406 14766 19458
rect 14030 19394 14082 19406
rect 15038 19394 15090 19406
rect 26126 19458 26178 19470
rect 26126 19394 26178 19406
rect 26350 19458 26402 19470
rect 26350 19394 26402 19406
rect 26910 19458 26962 19470
rect 26910 19394 26962 19406
rect 14478 19346 14530 19358
rect 25678 19346 25730 19358
rect 40014 19346 40066 19358
rect 22418 19294 22430 19346
rect 22482 19294 22494 19346
rect 24546 19294 24558 19346
rect 24610 19294 24622 19346
rect 26562 19294 26574 19346
rect 26626 19294 26638 19346
rect 14478 19282 14530 19294
rect 25678 19282 25730 19294
rect 40014 19282 40066 19294
rect 15150 19234 15202 19246
rect 26686 19234 26738 19246
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 15150 19170 15202 19182
rect 26686 19170 26738 19182
rect 27246 19234 27298 19246
rect 29374 19234 29426 19246
rect 30046 19234 30098 19246
rect 27794 19182 27806 19234
rect 27858 19182 27870 19234
rect 29698 19182 29710 19234
rect 29762 19182 29774 19234
rect 27246 19170 27298 19182
rect 29374 19170 29426 19182
rect 30046 19170 30098 19182
rect 30382 19234 30434 19246
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 30382 19170 30434 19182
rect 13806 19122 13858 19134
rect 13806 19058 13858 19070
rect 15038 19122 15090 19134
rect 24882 19070 24894 19122
rect 24946 19070 24958 19122
rect 15038 19058 15090 19070
rect 25230 19010 25282 19022
rect 25230 18946 25282 18958
rect 25566 19010 25618 19022
rect 25566 18946 25618 18958
rect 27358 19010 27410 19022
rect 27358 18946 27410 18958
rect 27470 19010 27522 19022
rect 27470 18946 27522 18958
rect 29150 19010 29202 19022
rect 29150 18946 29202 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 30158 19010 30210 19022
rect 30158 18946 30210 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 25342 18674 25394 18686
rect 25342 18610 25394 18622
rect 19294 18562 19346 18574
rect 24222 18562 24274 18574
rect 17714 18510 17726 18562
rect 17778 18510 17790 18562
rect 23874 18510 23886 18562
rect 23938 18510 23950 18562
rect 19294 18498 19346 18510
rect 24222 18498 24274 18510
rect 24334 18562 24386 18574
rect 24334 18498 24386 18510
rect 25230 18562 25282 18574
rect 25230 18498 25282 18510
rect 15150 18450 15202 18462
rect 23550 18450 23602 18462
rect 13906 18398 13918 18450
rect 13970 18398 13982 18450
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 17490 18398 17502 18450
rect 17554 18398 17566 18450
rect 19506 18398 19518 18450
rect 19570 18398 19582 18450
rect 27010 18398 27022 18450
rect 27074 18398 27086 18450
rect 27682 18398 27694 18450
rect 27746 18398 27758 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 15150 18386 15202 18398
rect 23550 18386 23602 18398
rect 25902 18338 25954 18350
rect 11778 18286 11790 18338
rect 11842 18286 11854 18338
rect 25902 18274 25954 18286
rect 26574 18338 26626 18350
rect 29810 18286 29822 18338
rect 29874 18286 29886 18338
rect 26574 18274 26626 18286
rect 24334 18226 24386 18238
rect 24334 18162 24386 18174
rect 25342 18226 25394 18238
rect 25342 18162 25394 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 19742 17890 19794 17902
rect 19742 17826 19794 17838
rect 19518 17778 19570 17790
rect 19518 17714 19570 17726
rect 15822 17666 15874 17678
rect 15698 17614 15710 17666
rect 15762 17614 15774 17666
rect 15822 17602 15874 17614
rect 15934 17666 15986 17678
rect 15934 17602 15986 17614
rect 16270 17666 16322 17678
rect 16270 17602 16322 17614
rect 16718 17666 16770 17678
rect 16718 17602 16770 17614
rect 16830 17666 16882 17678
rect 16830 17602 16882 17614
rect 17278 17666 17330 17678
rect 22642 17614 22654 17666
rect 22706 17614 22718 17666
rect 17278 17602 17330 17614
rect 23314 17502 23326 17554
rect 23378 17502 23390 17554
rect 15486 17442 15538 17454
rect 15486 17378 15538 17390
rect 16942 17442 16994 17454
rect 20066 17390 20078 17442
rect 20130 17390 20142 17442
rect 16942 17378 16994 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 18734 17106 18786 17118
rect 18734 17042 18786 17054
rect 18958 17106 19010 17118
rect 18958 17042 19010 17054
rect 22766 17106 22818 17118
rect 22766 17042 22818 17054
rect 22990 17106 23042 17118
rect 22990 17042 23042 17054
rect 23214 17106 23266 17118
rect 23214 17042 23266 17054
rect 17278 16994 17330 17006
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 17278 16930 17330 16942
rect 17502 16994 17554 17006
rect 17502 16930 17554 16942
rect 17614 16994 17666 17006
rect 17614 16930 17666 16942
rect 20414 16994 20466 17006
rect 26450 16942 26462 16994
rect 26514 16942 26526 16994
rect 20414 16930 20466 16942
rect 23662 16882 23714 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 20178 16830 20190 16882
rect 20242 16830 20254 16882
rect 23662 16818 23714 16830
rect 25342 16882 25394 16894
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 25342 16818 25394 16830
rect 18510 16770 18562 16782
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 18510 16706 18562 16718
rect 18846 16770 18898 16782
rect 18846 16706 18898 16718
rect 22878 16770 22930 16782
rect 22878 16706 22930 16718
rect 23886 16770 23938 16782
rect 28578 16718 28590 16770
rect 28642 16718 28654 16770
rect 23886 16706 23938 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 18286 16658 18338 16670
rect 24210 16606 24222 16658
rect 24274 16606 24286 16658
rect 18286 16594 18338 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 21310 16322 21362 16334
rect 21310 16258 21362 16270
rect 17054 16210 17106 16222
rect 13458 16158 13470 16210
rect 13522 16158 13534 16210
rect 15586 16158 15598 16210
rect 15650 16158 15662 16210
rect 17054 16146 17106 16158
rect 17502 16210 17554 16222
rect 26910 16210 26962 16222
rect 19058 16158 19070 16210
rect 19122 16158 19134 16210
rect 17502 16146 17554 16158
rect 26910 16146 26962 16158
rect 20190 16098 20242 16110
rect 16258 16046 16270 16098
rect 16322 16046 16334 16098
rect 19842 16046 19854 16098
rect 19906 16046 19918 16098
rect 20190 16034 20242 16046
rect 20638 16098 20690 16110
rect 20638 16034 20690 16046
rect 21422 16098 21474 16110
rect 23314 16046 23326 16098
rect 23378 16046 23390 16098
rect 21422 16034 21474 16046
rect 19294 15986 19346 15998
rect 20402 15934 20414 15986
rect 20466 15934 20478 15986
rect 24098 15934 24110 15986
rect 24162 15934 24174 15986
rect 19294 15922 19346 15934
rect 19070 15874 19122 15886
rect 21534 15874 21586 15886
rect 20178 15822 20190 15874
rect 20242 15822 20254 15874
rect 26338 15822 26350 15874
rect 26402 15822 26414 15874
rect 19070 15810 19122 15822
rect 21534 15810 21586 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 15710 15538 15762 15550
rect 15710 15474 15762 15486
rect 19294 15538 19346 15550
rect 19294 15474 19346 15486
rect 24110 15538 24162 15550
rect 24110 15474 24162 15486
rect 25230 15538 25282 15550
rect 25230 15474 25282 15486
rect 25902 15538 25954 15550
rect 25902 15474 25954 15486
rect 15598 15426 15650 15438
rect 19618 15374 19630 15426
rect 19682 15374 19694 15426
rect 21298 15374 21310 15426
rect 21362 15374 21374 15426
rect 25554 15374 25566 15426
rect 25618 15374 25630 15426
rect 26226 15374 26238 15426
rect 26290 15374 26302 15426
rect 15598 15362 15650 15374
rect 20514 15262 20526 15314
rect 20578 15262 20590 15314
rect 23874 15262 23886 15314
rect 23938 15262 23950 15314
rect 24558 15202 24610 15214
rect 23426 15150 23438 15202
rect 23490 15150 23502 15202
rect 24558 15138 24610 15150
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19966 14642 20018 14654
rect 17378 14590 17390 14642
rect 17442 14590 17454 14642
rect 19506 14590 19518 14642
rect 19570 14590 19582 14642
rect 19966 14578 20018 14590
rect 16594 14478 16606 14530
rect 16658 14478 16670 14530
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 22318 13970 22370 13982
rect 22318 13906 22370 13918
rect 19730 13806 19742 13858
rect 19794 13806 19806 13858
rect 18946 13694 18958 13746
rect 19010 13694 19022 13746
rect 21858 13582 21870 13634
rect 21922 13582 21934 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 18062 5234 18114 5246
rect 18062 5170 18114 5182
rect 17042 5070 17054 5122
rect 17106 5070 17118 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 19730 4286 19742 4338
rect 19794 4286 19806 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 20750 4114 20802 4126
rect 20750 4050 20802 4062
rect 26798 4114 26850 4126
rect 26798 4050 26850 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 22430 3666 22482 3678
rect 18834 3614 18846 3666
rect 18898 3614 18910 3666
rect 22430 3602 22482 3614
rect 24782 3666 24834 3678
rect 24782 3602 24834 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 21746 3502 21758 3554
rect 21810 3502 21822 3554
rect 27010 3502 27022 3554
rect 27074 3502 27086 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19518 38222 19570 38274
rect 22094 38222 22146 38274
rect 17614 37998 17666 38050
rect 21310 37998 21362 38050
rect 16942 37886 16994 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18510 37438 18562 37490
rect 21422 37438 21474 37490
rect 17502 37214 17554 37266
rect 20862 37214 20914 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 40238 36318 40290 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 20750 27134 20802 27186
rect 17950 27022 18002 27074
rect 21646 27022 21698 27074
rect 18622 26910 18674 26962
rect 21310 26910 21362 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17390 26350 17442 26402
rect 13918 26238 13970 26290
rect 26574 26238 26626 26290
rect 37662 26238 37714 26290
rect 14702 26126 14754 26178
rect 16830 26126 16882 26178
rect 17950 26126 18002 26178
rect 20974 26126 21026 26178
rect 24334 26126 24386 26178
rect 26238 26126 26290 26178
rect 27358 26126 27410 26178
rect 29486 26126 29538 26178
rect 39902 26126 39954 26178
rect 17502 26014 17554 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 27358 25678 27410 25730
rect 1934 25566 1986 25618
rect 16606 25566 16658 25618
rect 22542 25566 22594 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 13470 25454 13522 25506
rect 19406 25454 19458 25506
rect 25342 25454 25394 25506
rect 27470 25454 27522 25506
rect 29262 25454 29314 25506
rect 37662 25454 37714 25506
rect 13806 25342 13858 25394
rect 18734 25342 18786 25394
rect 24670 25342 24722 25394
rect 27918 25342 27970 25394
rect 28030 25342 28082 25394
rect 13694 25230 13746 25282
rect 19966 25230 20018 25282
rect 25902 25230 25954 25282
rect 26350 25230 26402 25282
rect 27358 25230 27410 25282
rect 27694 25230 27746 25282
rect 29486 25230 29538 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15262 24894 15314 24946
rect 15374 24894 15426 24946
rect 17614 24894 17666 24946
rect 17726 24894 17778 24946
rect 18846 24894 18898 24946
rect 19294 24894 19346 24946
rect 20414 24894 20466 24946
rect 24782 24894 24834 24946
rect 13918 24782 13970 24834
rect 18958 24782 19010 24834
rect 24558 24782 24610 24834
rect 14702 24670 14754 24722
rect 15038 24670 15090 24722
rect 15486 24670 15538 24722
rect 15710 24670 15762 24722
rect 17502 24670 17554 24722
rect 17838 24670 17890 24722
rect 17950 24670 18002 24722
rect 19518 24670 19570 24722
rect 19742 24670 19794 24722
rect 20078 24670 20130 24722
rect 20302 24670 20354 24722
rect 20638 24670 20690 24722
rect 20974 24670 21026 24722
rect 21198 24670 21250 24722
rect 24446 24670 24498 24722
rect 25566 24670 25618 24722
rect 37662 24670 37714 24722
rect 11790 24558 11842 24610
rect 21982 24558 22034 24610
rect 24110 24558 24162 24610
rect 26350 24558 26402 24610
rect 28478 24558 28530 24610
rect 18846 24446 18898 24498
rect 19630 24446 19682 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 13470 24110 13522 24162
rect 27022 24110 27074 24162
rect 1934 23998 1986 24050
rect 18622 23998 18674 24050
rect 23550 23998 23602 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 13806 23886 13858 23938
rect 18734 23886 18786 23938
rect 18958 23886 19010 23938
rect 19182 23886 19234 23938
rect 19406 23886 19458 23938
rect 22654 23886 22706 23938
rect 27134 23886 27186 23938
rect 28142 23886 28194 23938
rect 28478 23886 28530 23938
rect 29374 23886 29426 23938
rect 37662 23886 37714 23938
rect 18510 23774 18562 23826
rect 27022 23774 27074 23826
rect 28366 23774 28418 23826
rect 13582 23662 13634 23714
rect 14926 23662 14978 23714
rect 29038 23662 29090 23714
rect 29262 23662 29314 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 14926 23326 14978 23378
rect 15150 23326 15202 23378
rect 15934 23326 15986 23378
rect 21758 23326 21810 23378
rect 21870 23326 21922 23378
rect 23102 23326 23154 23378
rect 26798 23326 26850 23378
rect 13694 23214 13746 23266
rect 15486 23214 15538 23266
rect 21086 23214 21138 23266
rect 21982 23214 22034 23266
rect 22766 23214 22818 23266
rect 14478 23102 14530 23154
rect 15038 23102 15090 23154
rect 15262 23102 15314 23154
rect 20414 23102 20466 23154
rect 20638 23102 20690 23154
rect 21310 23102 21362 23154
rect 22430 23102 22482 23154
rect 23662 23102 23714 23154
rect 24110 23102 24162 23154
rect 27134 23102 27186 23154
rect 11566 22990 11618 23042
rect 19742 22990 19794 23042
rect 24222 22990 24274 23042
rect 27918 22990 27970 23042
rect 30046 22990 30098 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 15486 22542 15538 22594
rect 18734 22542 18786 22594
rect 21310 22542 21362 22594
rect 21646 22542 21698 22594
rect 22318 22542 22370 22594
rect 27918 22542 27970 22594
rect 1934 22430 1986 22482
rect 21870 22430 21922 22482
rect 24558 22430 24610 22482
rect 4286 22318 4338 22370
rect 14030 22318 14082 22370
rect 14254 22318 14306 22370
rect 15486 22318 15538 22370
rect 17614 22318 17666 22370
rect 17838 22318 17890 22370
rect 24334 22318 24386 22370
rect 28030 22318 28082 22370
rect 12686 22206 12738 22258
rect 12910 22206 12962 22258
rect 14142 22206 14194 22258
rect 14590 22206 14642 22258
rect 15150 22206 15202 22258
rect 16942 22206 16994 22258
rect 17278 22206 17330 22258
rect 18062 22206 18114 22258
rect 18398 22206 18450 22258
rect 18846 22206 18898 22258
rect 22206 22206 22258 22258
rect 23662 22206 23714 22258
rect 24110 22206 24162 22258
rect 12798 22094 12850 22146
rect 18174 22094 18226 22146
rect 18622 22094 18674 22146
rect 22318 22094 22370 22146
rect 27918 22094 27970 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 16606 21758 16658 21810
rect 17726 21758 17778 21810
rect 19630 21758 19682 21810
rect 22766 21758 22818 21810
rect 13134 21646 13186 21698
rect 17390 21646 17442 21698
rect 19182 21646 19234 21698
rect 19742 21646 19794 21698
rect 20638 21646 20690 21698
rect 21534 21646 21586 21698
rect 22206 21646 22258 21698
rect 22990 21646 23042 21698
rect 23774 21646 23826 21698
rect 24222 21646 24274 21698
rect 24670 21646 24722 21698
rect 25230 21646 25282 21698
rect 27806 21646 27858 21698
rect 13918 21534 13970 21586
rect 14366 21534 14418 21586
rect 16830 21534 16882 21586
rect 18398 21534 18450 21586
rect 18734 21534 18786 21586
rect 19966 21534 20018 21586
rect 20190 21534 20242 21586
rect 21758 21534 21810 21586
rect 22430 21534 22482 21586
rect 23102 21534 23154 21586
rect 24446 21534 24498 21586
rect 25566 21534 25618 21586
rect 27582 21534 27634 21586
rect 27918 21534 27970 21586
rect 37662 21534 37714 21586
rect 11006 21422 11058 21474
rect 19182 21422 19234 21474
rect 16494 21310 16546 21362
rect 20526 21310 20578 21362
rect 40014 21310 40066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 19406 20974 19458 21026
rect 1934 20862 1986 20914
rect 16046 20862 16098 20914
rect 16382 20862 16434 20914
rect 17950 20862 18002 20914
rect 23550 20862 23602 20914
rect 4174 20750 4226 20802
rect 14926 20750 14978 20802
rect 15262 20750 15314 20802
rect 16718 20750 16770 20802
rect 19070 20750 19122 20802
rect 19966 20750 20018 20802
rect 21310 20750 21362 20802
rect 15486 20638 15538 20690
rect 16158 20638 16210 20690
rect 17166 20638 17218 20690
rect 19742 20638 19794 20690
rect 20414 20638 20466 20690
rect 20526 20638 20578 20690
rect 15598 20526 15650 20578
rect 16830 20526 16882 20578
rect 16942 20526 16994 20578
rect 17838 20526 17890 20578
rect 18062 20526 18114 20578
rect 18286 20526 18338 20578
rect 19294 20526 19346 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14590 20190 14642 20242
rect 18622 20190 18674 20242
rect 18958 20190 19010 20242
rect 22430 20190 22482 20242
rect 23102 20190 23154 20242
rect 15486 20078 15538 20130
rect 16046 20078 16098 20130
rect 19406 20078 19458 20130
rect 19630 20078 19682 20130
rect 19966 20078 20018 20130
rect 21086 20078 21138 20130
rect 21982 20078 22034 20130
rect 24446 20078 24498 20130
rect 25342 20078 25394 20130
rect 28926 20078 28978 20130
rect 29598 20078 29650 20130
rect 29710 20078 29762 20130
rect 4286 19966 4338 20018
rect 14254 19966 14306 20018
rect 14814 19966 14866 20018
rect 15262 19966 15314 20018
rect 15710 19966 15762 20018
rect 19294 19966 19346 20018
rect 19854 19966 19906 20018
rect 21422 19966 21474 20018
rect 21534 19966 21586 20018
rect 21870 19966 21922 20018
rect 22206 19966 22258 20018
rect 22766 19966 22818 20018
rect 23326 19966 23378 20018
rect 24222 19966 24274 20018
rect 25678 19966 25730 20018
rect 29150 19966 29202 20018
rect 11342 19854 11394 19906
rect 13470 19854 13522 19906
rect 14702 19854 14754 19906
rect 15598 19854 15650 19906
rect 26462 19854 26514 19906
rect 28590 19854 28642 19906
rect 1934 19742 1986 19794
rect 19966 19742 20018 19794
rect 29710 19742 29762 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 13694 19406 13746 19458
rect 14030 19406 14082 19458
rect 14254 19406 14306 19458
rect 14702 19406 14754 19458
rect 15038 19406 15090 19458
rect 26126 19406 26178 19458
rect 26350 19406 26402 19458
rect 26910 19406 26962 19458
rect 14478 19294 14530 19346
rect 22430 19294 22482 19346
rect 24558 19294 24610 19346
rect 25678 19294 25730 19346
rect 26574 19294 26626 19346
rect 40014 19294 40066 19346
rect 15150 19182 15202 19234
rect 21758 19182 21810 19234
rect 26686 19182 26738 19234
rect 27246 19182 27298 19234
rect 27806 19182 27858 19234
rect 29374 19182 29426 19234
rect 29710 19182 29762 19234
rect 30046 19182 30098 19234
rect 30382 19182 30434 19234
rect 37662 19182 37714 19234
rect 13806 19070 13858 19122
rect 15038 19070 15090 19122
rect 24894 19070 24946 19122
rect 25230 18958 25282 19010
rect 25566 18958 25618 19010
rect 27358 18958 27410 19010
rect 27470 18958 27522 19010
rect 29150 18958 29202 19010
rect 29262 18958 29314 19010
rect 30158 18958 30210 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 25342 18622 25394 18674
rect 17726 18510 17778 18562
rect 19294 18510 19346 18562
rect 23886 18510 23938 18562
rect 24222 18510 24274 18562
rect 24334 18510 24386 18562
rect 25230 18510 25282 18562
rect 13918 18398 13970 18450
rect 14590 18398 14642 18450
rect 15150 18398 15202 18450
rect 17502 18398 17554 18450
rect 19518 18398 19570 18450
rect 23550 18398 23602 18450
rect 27022 18398 27074 18450
rect 27694 18398 27746 18450
rect 37662 18398 37714 18450
rect 11790 18286 11842 18338
rect 25902 18286 25954 18338
rect 26574 18286 26626 18338
rect 29822 18286 29874 18338
rect 24334 18174 24386 18226
rect 25342 18174 25394 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 19742 17838 19794 17890
rect 19518 17726 19570 17778
rect 15710 17614 15762 17666
rect 15822 17614 15874 17666
rect 15934 17614 15986 17666
rect 16270 17614 16322 17666
rect 16718 17614 16770 17666
rect 16830 17614 16882 17666
rect 17278 17614 17330 17666
rect 22654 17614 22706 17666
rect 23326 17502 23378 17554
rect 15486 17390 15538 17442
rect 16942 17390 16994 17442
rect 20078 17390 20130 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 18734 17054 18786 17106
rect 18958 17054 19010 17106
rect 22766 17054 22818 17106
rect 22990 17054 23042 17106
rect 23214 17054 23266 17106
rect 14702 16942 14754 16994
rect 17278 16942 17330 16994
rect 17502 16942 17554 16994
rect 17614 16942 17666 16994
rect 20414 16942 20466 16994
rect 26462 16942 26514 16994
rect 4286 16830 4338 16882
rect 14030 16830 14082 16882
rect 20190 16830 20242 16882
rect 23662 16830 23714 16882
rect 25342 16830 25394 16882
rect 25790 16830 25842 16882
rect 16830 16718 16882 16770
rect 18510 16718 18562 16770
rect 18846 16718 18898 16770
rect 22878 16718 22930 16770
rect 23886 16718 23938 16770
rect 28590 16718 28642 16770
rect 1934 16606 1986 16658
rect 18286 16606 18338 16658
rect 24222 16606 24274 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 21310 16270 21362 16322
rect 13470 16158 13522 16210
rect 15598 16158 15650 16210
rect 17054 16158 17106 16210
rect 17502 16158 17554 16210
rect 19070 16158 19122 16210
rect 26910 16158 26962 16210
rect 16270 16046 16322 16098
rect 19854 16046 19906 16098
rect 20190 16046 20242 16098
rect 20638 16046 20690 16098
rect 21422 16046 21474 16098
rect 23326 16046 23378 16098
rect 19294 15934 19346 15986
rect 20414 15934 20466 15986
rect 24110 15934 24162 15986
rect 19070 15822 19122 15874
rect 20190 15822 20242 15874
rect 21534 15822 21586 15874
rect 26350 15822 26402 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 15710 15486 15762 15538
rect 19294 15486 19346 15538
rect 24110 15486 24162 15538
rect 25230 15486 25282 15538
rect 25902 15486 25954 15538
rect 15598 15374 15650 15426
rect 19630 15374 19682 15426
rect 21310 15374 21362 15426
rect 25566 15374 25618 15426
rect 26238 15374 26290 15426
rect 20526 15262 20578 15314
rect 23886 15262 23938 15314
rect 23438 15150 23490 15202
rect 24558 15150 24610 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 17390 14590 17442 14642
rect 19518 14590 19570 14642
rect 19966 14590 20018 14642
rect 16606 14478 16658 14530
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 22318 13918 22370 13970
rect 19742 13806 19794 13858
rect 18958 13694 19010 13746
rect 21870 13582 21922 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 18062 5182 18114 5234
rect 17054 5070 17106 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19742 4286 19794 4338
rect 25790 4286 25842 4338
rect 20750 4062 20802 4114
rect 26798 4062 26850 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18846 3614 18898 3666
rect 22430 3614 22482 3666
rect 24782 3614 24834 3666
rect 29374 3614 29426 3666
rect 19742 3502 19794 3554
rect 21758 3502 21810 3554
rect 27022 3502 27074 3554
rect 28590 3502 28642 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16128 41200 16240 42000
rect 17472 41200 17584 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 20832 41200 20944 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 16156 37940 16212 41200
rect 16156 37874 16212 37884
rect 16940 37940 16996 37950
rect 16940 37846 16996 37884
rect 17500 37492 17556 41200
rect 19516 38274 19572 41200
rect 19516 38222 19518 38274
rect 19570 38222 19572 38274
rect 19516 38210 19572 38222
rect 17500 37426 17556 37436
rect 17612 38050 17668 38062
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 17500 37266 17556 37278
rect 17500 37214 17502 37266
rect 17554 37214 17556 37266
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 17500 31948 17556 37214
rect 17388 31892 17556 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 17388 26404 17444 31892
rect 16828 26402 17444 26404
rect 16828 26350 17390 26402
rect 17442 26350 17444 26402
rect 16828 26348 17444 26350
rect 4172 26292 4228 26302
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22484 1988 22494
rect 1932 22390 1988 22428
rect 4172 21028 4228 26236
rect 13916 26290 13972 26302
rect 13916 26238 13918 26290
rect 13970 26238 13972 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 11788 25508 11844 25518
rect 11788 24948 11844 25452
rect 11788 24610 11844 24892
rect 11788 24558 11790 24610
rect 11842 24558 11844 24610
rect 11788 24546 11844 24558
rect 13468 25506 13524 25518
rect 13468 25454 13470 25506
rect 13522 25454 13524 25506
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 12684 24276 12740 24286
rect 4284 23938 4340 23950
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23044 4340 23886
rect 4284 22978 4340 22988
rect 11564 23156 11620 23166
rect 11564 23042 11620 23100
rect 11564 22990 11566 23042
rect 11618 22990 11620 23042
rect 11564 22978 11620 22990
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22372 4340 22382
rect 4284 22278 4340 22316
rect 11004 22372 11060 22382
rect 11004 21474 11060 22316
rect 12684 22258 12740 24220
rect 13468 24276 13524 25454
rect 13804 25394 13860 25406
rect 13804 25342 13806 25394
rect 13858 25342 13860 25394
rect 13692 25282 13748 25294
rect 13692 25230 13694 25282
rect 13746 25230 13748 25282
rect 13692 24948 13748 25230
rect 13804 25172 13860 25342
rect 13916 25284 13972 26238
rect 14700 26180 14756 26190
rect 14700 26178 14868 26180
rect 14700 26126 14702 26178
rect 14754 26126 14868 26178
rect 14700 26124 14868 26126
rect 14700 26114 14756 26124
rect 13916 25218 13972 25228
rect 14700 25284 14756 25294
rect 13804 25106 13860 25116
rect 13692 24892 13972 24948
rect 13916 24834 13972 24892
rect 13916 24782 13918 24834
rect 13970 24782 13972 24834
rect 13916 24770 13972 24782
rect 14700 24724 14756 25228
rect 14812 25060 14868 26124
rect 16828 26178 16884 26348
rect 17388 26338 17444 26348
rect 16828 26126 16830 26178
rect 16882 26126 16884 26178
rect 16828 26114 16884 26126
rect 17500 26066 17556 26078
rect 17500 26014 17502 26066
rect 17554 26014 17556 26066
rect 16604 25620 16660 25630
rect 16604 25526 16660 25564
rect 14812 24994 14868 25004
rect 15372 25172 15428 25182
rect 15260 24948 15316 24958
rect 15260 24854 15316 24892
rect 15372 24946 15428 25116
rect 15372 24894 15374 24946
rect 15426 24894 15428 24946
rect 15372 24882 15428 24894
rect 17500 24948 17556 26014
rect 17612 25620 17668 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18508 37492 18564 37502
rect 18508 37398 18564 37436
rect 20188 37492 20244 41200
rect 20860 38276 20916 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 20860 38210 20916 38220
rect 22092 38276 22148 38286
rect 22092 38182 22148 38220
rect 20188 37426 20244 37436
rect 21308 38050 21364 38062
rect 21308 37998 21310 38050
rect 21362 37998 21364 38050
rect 20860 37268 20916 37278
rect 20860 37174 20916 37212
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20748 27186 20804 27198
rect 20748 27134 20750 27186
rect 20802 27134 20804 27186
rect 17612 25554 17668 25564
rect 17948 27074 18004 27086
rect 17948 27022 17950 27074
rect 18002 27022 18004 27074
rect 17948 26178 18004 27022
rect 18620 26962 18676 26974
rect 18620 26910 18622 26962
rect 18674 26910 18676 26962
rect 18620 26908 18676 26910
rect 20748 26908 20804 27134
rect 21308 26962 21364 37998
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 18620 26852 19348 26908
rect 17948 26126 17950 26178
rect 18002 26126 18004 26178
rect 17948 25284 18004 26126
rect 18844 25620 18900 25630
rect 18732 25396 18788 25406
rect 17948 25218 18004 25228
rect 18620 25394 18788 25396
rect 18620 25342 18734 25394
rect 18786 25342 18788 25394
rect 18620 25340 18788 25342
rect 17724 25060 17780 25070
rect 17612 24948 17668 24958
rect 17500 24946 17668 24948
rect 17500 24894 17614 24946
rect 17666 24894 17668 24946
rect 17500 24892 17668 24894
rect 17612 24882 17668 24892
rect 17724 24946 17780 25004
rect 17724 24894 17726 24946
rect 17778 24894 17780 24946
rect 17724 24882 17780 24894
rect 15036 24724 15092 24734
rect 14700 24722 14868 24724
rect 14700 24670 14702 24722
rect 14754 24670 14868 24722
rect 14700 24668 14868 24670
rect 14700 24658 14756 24668
rect 13468 24162 13524 24220
rect 13468 24110 13470 24162
rect 13522 24110 13524 24162
rect 13468 24098 13524 24110
rect 13804 23940 13860 23950
rect 13804 23846 13860 23884
rect 13580 23714 13636 23726
rect 13580 23662 13582 23714
rect 13634 23662 13636 23714
rect 13580 23268 13636 23662
rect 14812 23716 14868 24668
rect 15036 24630 15092 24668
rect 15484 24722 15540 24734
rect 15484 24670 15486 24722
rect 15538 24670 15540 24722
rect 14924 23940 14980 23950
rect 14980 23884 15092 23940
rect 14924 23874 14980 23884
rect 14924 23716 14980 23726
rect 14812 23714 14980 23716
rect 14812 23662 14926 23714
rect 14978 23662 14980 23714
rect 14812 23660 14980 23662
rect 14028 23604 14084 23614
rect 13692 23268 13748 23278
rect 13580 23266 13748 23268
rect 13580 23214 13694 23266
rect 13746 23214 13748 23266
rect 13580 23212 13748 23214
rect 13692 23202 13748 23212
rect 14028 22370 14084 23548
rect 14812 23380 14868 23660
rect 14924 23650 14980 23660
rect 14476 23156 14532 23166
rect 14812 23156 14868 23324
rect 14924 23492 14980 23502
rect 14924 23378 14980 23436
rect 14924 23326 14926 23378
rect 14978 23326 14980 23378
rect 14924 23314 14980 23326
rect 15036 23380 15092 23884
rect 15148 23380 15204 23390
rect 15036 23378 15204 23380
rect 15036 23326 15150 23378
rect 15202 23326 15204 23378
rect 15036 23324 15204 23326
rect 15148 23314 15204 23324
rect 15484 23266 15540 24670
rect 15708 24722 15764 24734
rect 15708 24670 15710 24722
rect 15762 24670 15764 24722
rect 15708 23716 15764 24670
rect 17500 24724 17556 24734
rect 15708 23650 15764 23660
rect 17388 23716 17444 23726
rect 15932 23380 15988 23390
rect 15932 23286 15988 23324
rect 15484 23214 15486 23266
rect 15538 23214 15540 23266
rect 14476 23154 14868 23156
rect 14476 23102 14478 23154
rect 14530 23102 14868 23154
rect 14476 23100 14868 23102
rect 15036 23156 15092 23166
rect 14028 22318 14030 22370
rect 14082 22318 14084 22370
rect 14028 22306 14084 22318
rect 14252 22372 14308 22382
rect 14252 22278 14308 22316
rect 12684 22206 12686 22258
rect 12738 22206 12740 22258
rect 12684 22194 12740 22206
rect 12908 22260 12964 22270
rect 12908 22166 12964 22204
rect 14140 22260 14196 22270
rect 14140 22166 14196 22204
rect 12796 22146 12852 22158
rect 12796 22094 12798 22146
rect 12850 22094 12852 22146
rect 12796 21812 12852 22094
rect 12796 21756 13188 21812
rect 13132 21698 13188 21756
rect 13132 21646 13134 21698
rect 13186 21646 13188 21698
rect 13132 21634 13188 21646
rect 13916 21588 13972 21598
rect 14364 21588 14420 21598
rect 14476 21588 14532 23100
rect 15036 23062 15092 23100
rect 15260 23156 15316 23166
rect 15260 23062 15316 23100
rect 15484 22594 15540 23214
rect 15484 22542 15486 22594
rect 15538 22542 15540 22594
rect 15484 22530 15540 22542
rect 16604 23156 16660 23166
rect 15484 22370 15540 22382
rect 15484 22318 15486 22370
rect 15538 22318 15540 22370
rect 13916 21586 14532 21588
rect 13916 21534 13918 21586
rect 13970 21534 14366 21586
rect 14418 21534 14532 21586
rect 13916 21532 14532 21534
rect 14588 22258 14644 22270
rect 14588 22206 14590 22258
rect 14642 22206 14644 22258
rect 13916 21522 13972 21532
rect 14364 21522 14420 21532
rect 11004 21422 11006 21474
rect 11058 21422 11060 21474
rect 11004 21410 11060 21422
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 14588 21140 14644 22206
rect 14588 21074 14644 21084
rect 15148 22258 15204 22270
rect 15148 22206 15150 22258
rect 15202 22206 15204 22258
rect 4172 20962 4228 20972
rect 1932 20914 1988 20926
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20244 1988 20862
rect 1932 20178 1988 20188
rect 4172 20802 4228 20814
rect 4172 20750 4174 20802
rect 4226 20750 4228 20802
rect 4172 19908 4228 20750
rect 14924 20802 14980 20814
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 13804 20692 13860 20702
rect 11788 20132 11844 20142
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 11340 20020 11396 20030
rect 4172 19842 4228 19852
rect 11340 19906 11396 19964
rect 11340 19854 11342 19906
rect 11394 19854 11396 19906
rect 11340 19842 11396 19854
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 11788 19124 11844 20076
rect 13468 19908 13524 19918
rect 13468 19906 13748 19908
rect 13468 19854 13470 19906
rect 13522 19854 13748 19906
rect 13468 19852 13748 19854
rect 13468 19842 13524 19852
rect 13692 19458 13748 19852
rect 13692 19406 13694 19458
rect 13746 19406 13748 19458
rect 13692 19394 13748 19406
rect 11788 18338 11844 19068
rect 13804 19122 13860 20636
rect 14924 20692 14980 20750
rect 15148 20804 15204 22206
rect 15484 22260 15540 22318
rect 16604 22372 16660 23100
rect 15260 20804 15316 20814
rect 15148 20748 15260 20804
rect 15260 20710 15316 20748
rect 14924 20626 14980 20636
rect 15484 20690 15540 22204
rect 16156 22260 16212 22270
rect 15484 20638 15486 20690
rect 15538 20638 15540 20690
rect 15484 20626 15540 20638
rect 15932 21140 15988 21150
rect 15932 20916 15988 21084
rect 16044 20916 16100 20926
rect 15932 20914 16100 20916
rect 15932 20862 16046 20914
rect 16098 20862 16100 20914
rect 15932 20860 16100 20862
rect 15596 20578 15652 20590
rect 15596 20526 15598 20578
rect 15650 20526 15652 20578
rect 14588 20244 14644 20254
rect 14588 20150 14644 20188
rect 15260 20132 15316 20142
rect 14252 20020 14308 20030
rect 14812 20020 14868 20030
rect 14252 20018 14532 20020
rect 14252 19966 14254 20018
rect 14306 19966 14532 20018
rect 14252 19964 14532 19966
rect 14252 19954 14308 19964
rect 13804 19070 13806 19122
rect 13858 19070 13860 19122
rect 13804 19058 13860 19070
rect 13916 19908 13972 19918
rect 13916 18450 13972 19852
rect 14028 19460 14084 19470
rect 14252 19460 14308 19470
rect 14028 19458 14308 19460
rect 14028 19406 14030 19458
rect 14082 19406 14254 19458
rect 14306 19406 14308 19458
rect 14028 19404 14308 19406
rect 14028 19394 14084 19404
rect 14252 19394 14308 19404
rect 14476 19346 14532 19964
rect 14812 19926 14868 19964
rect 15036 20020 15092 20030
rect 14700 19906 14756 19918
rect 14700 19854 14702 19906
rect 14754 19854 14756 19906
rect 14700 19458 14756 19854
rect 14700 19406 14702 19458
rect 14754 19406 14756 19458
rect 14700 19394 14756 19406
rect 15036 19458 15092 19964
rect 15260 20018 15316 20076
rect 15484 20132 15540 20142
rect 15596 20132 15652 20526
rect 15484 20130 15652 20132
rect 15484 20078 15486 20130
rect 15538 20078 15652 20130
rect 15484 20076 15652 20078
rect 15484 20066 15540 20076
rect 15260 19966 15262 20018
rect 15314 19966 15316 20018
rect 15260 19954 15316 19966
rect 15708 20020 15764 20030
rect 15708 19926 15764 19964
rect 15596 19908 15652 19918
rect 15596 19814 15652 19852
rect 15932 19796 15988 20860
rect 16044 20850 16100 20860
rect 16156 20690 16212 22204
rect 16604 21810 16660 22316
rect 16940 22260 16996 22270
rect 16940 22166 16996 22204
rect 17276 22258 17332 22270
rect 17276 22206 17278 22258
rect 17330 22206 17332 22258
rect 16604 21758 16606 21810
rect 16658 21758 16660 21810
rect 16604 21746 16660 21758
rect 17276 21700 17332 22206
rect 16828 21588 16884 21598
rect 17164 21588 17220 21598
rect 16828 21586 17164 21588
rect 16828 21534 16830 21586
rect 16882 21534 17164 21586
rect 16828 21532 17164 21534
rect 16828 21522 16884 21532
rect 16492 21362 16548 21374
rect 16492 21310 16494 21362
rect 16546 21310 16548 21362
rect 16380 20916 16436 20926
rect 16492 20916 16548 21310
rect 16380 20914 16492 20916
rect 16380 20862 16382 20914
rect 16434 20862 16492 20914
rect 16380 20860 16492 20862
rect 16380 20850 16436 20860
rect 16492 20850 16548 20860
rect 16716 21140 16772 21150
rect 16716 20804 16772 21084
rect 16716 20710 16772 20748
rect 16156 20638 16158 20690
rect 16210 20638 16212 20690
rect 16156 20626 16212 20638
rect 17164 20690 17220 21532
rect 17164 20638 17166 20690
rect 17218 20638 17220 20690
rect 17164 20626 17220 20638
rect 16828 20578 16884 20590
rect 16828 20526 16830 20578
rect 16882 20526 16884 20578
rect 16044 20244 16100 20254
rect 16044 20130 16100 20188
rect 16044 20078 16046 20130
rect 16098 20078 16100 20130
rect 16044 20066 16100 20078
rect 16828 20132 16884 20526
rect 16940 20580 16996 20590
rect 16940 20578 17108 20580
rect 16940 20526 16942 20578
rect 16994 20526 17108 20578
rect 16940 20524 17108 20526
rect 16940 20514 16996 20524
rect 17052 20468 17108 20524
rect 17276 20468 17332 21644
rect 17388 21698 17444 23660
rect 17500 23604 17556 24668
rect 17836 24724 17892 24734
rect 17836 24630 17892 24668
rect 17948 24722 18004 24734
rect 17948 24670 17950 24722
rect 18002 24670 18004 24722
rect 17500 23538 17556 23548
rect 17612 22372 17668 22382
rect 17612 22278 17668 22316
rect 17836 22372 17892 22382
rect 17836 22278 17892 22316
rect 17948 21924 18004 24670
rect 18620 24050 18676 25340
rect 18732 25330 18788 25340
rect 18844 24946 18900 25564
rect 18844 24894 18846 24946
rect 18898 24894 18900 24946
rect 18844 24882 18900 24894
rect 19292 24946 19348 26852
rect 20412 26852 21252 26908
rect 21308 26898 21364 26910
rect 21644 37268 21700 37278
rect 21644 27074 21700 37212
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 40236 36372 40292 36382
rect 40236 36278 40292 36316
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 21644 27022 21646 27074
rect 21698 27022 21700 27074
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19404 25506 19460 25518
rect 19404 25454 19406 25506
rect 19458 25454 19460 25506
rect 19404 25284 19460 25454
rect 19404 25218 19460 25228
rect 19964 25284 20020 25322
rect 19964 25218 20020 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19292 24894 19294 24946
rect 19346 24894 19348 24946
rect 19292 24882 19348 24894
rect 20412 24946 20468 26852
rect 21196 26740 21252 26852
rect 21644 26740 21700 27022
rect 21196 26684 21700 26740
rect 26572 26290 26628 26302
rect 26572 26238 26574 26290
rect 26626 26238 26628 26290
rect 20972 26178 21028 26190
rect 20972 26126 20974 26178
rect 21026 26126 21028 26178
rect 20972 25284 21028 26126
rect 24332 26178 24388 26190
rect 24332 26126 24334 26178
rect 24386 26126 24388 26178
rect 22540 25618 22596 25630
rect 22540 25566 22542 25618
rect 22594 25566 22596 25618
rect 21028 25228 21252 25284
rect 20972 25218 21028 25228
rect 20412 24894 20414 24946
rect 20466 24894 20468 24946
rect 20412 24882 20468 24894
rect 18956 24836 19012 24846
rect 18956 24742 19012 24780
rect 20972 24836 21028 24846
rect 18732 24724 18788 24734
rect 18732 24164 18788 24668
rect 19516 24722 19572 24734
rect 19516 24670 19518 24722
rect 19570 24670 19572 24722
rect 18844 24500 18900 24510
rect 18844 24498 19460 24500
rect 18844 24446 18846 24498
rect 18898 24446 19460 24498
rect 18844 24444 19460 24446
rect 18844 24434 18900 24444
rect 18732 24108 18900 24164
rect 18620 23998 18622 24050
rect 18674 23998 18676 24050
rect 18620 23986 18676 23998
rect 18732 23938 18788 23950
rect 18732 23886 18734 23938
rect 18786 23886 18788 23938
rect 18508 23826 18564 23838
rect 18508 23774 18510 23826
rect 18562 23774 18564 23826
rect 18060 22260 18116 22270
rect 18060 22166 18116 22204
rect 18396 22260 18452 22270
rect 18508 22260 18564 23774
rect 18732 23716 18788 23886
rect 18732 23650 18788 23660
rect 18732 22596 18788 22606
rect 18844 22596 18900 24108
rect 18956 23938 19012 23950
rect 18956 23886 18958 23938
rect 19010 23886 19012 23938
rect 18956 23044 19012 23886
rect 19180 23940 19236 23950
rect 19180 23846 19236 23884
rect 19404 23938 19460 24444
rect 19516 24276 19572 24670
rect 19740 24724 19796 24734
rect 19740 24630 19796 24668
rect 20076 24724 20132 24734
rect 20300 24724 20356 24734
rect 20076 24722 20356 24724
rect 20076 24670 20078 24722
rect 20130 24670 20302 24722
rect 20354 24670 20356 24722
rect 20076 24668 20356 24670
rect 20076 24658 20132 24668
rect 20300 24658 20356 24668
rect 20636 24722 20692 24734
rect 20636 24670 20638 24722
rect 20690 24670 20692 24722
rect 19516 24210 19572 24220
rect 19628 24498 19684 24510
rect 19628 24446 19630 24498
rect 19682 24446 19684 24498
rect 19404 23886 19406 23938
rect 19458 23886 19460 23938
rect 19404 23874 19460 23886
rect 19516 23940 19572 23950
rect 18956 22978 19012 22988
rect 19180 23604 19236 23614
rect 18732 22594 18900 22596
rect 18732 22542 18734 22594
rect 18786 22542 18900 22594
rect 18732 22540 18900 22542
rect 18732 22530 18788 22540
rect 18844 22260 18900 22270
rect 18452 22204 18564 22260
rect 18732 22258 18900 22260
rect 18732 22206 18846 22258
rect 18898 22206 18900 22258
rect 18732 22204 18900 22206
rect 18396 22166 18452 22204
rect 18172 22148 18228 22158
rect 18172 22054 18228 22092
rect 18620 22146 18676 22158
rect 18620 22094 18622 22146
rect 18674 22094 18676 22146
rect 17836 21868 18004 21924
rect 17724 21812 17780 21822
rect 17724 21718 17780 21756
rect 17388 21646 17390 21698
rect 17442 21646 17444 21698
rect 17388 20692 17444 21646
rect 17836 20916 17892 21868
rect 18396 21812 18452 21822
rect 18396 21586 18452 21756
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 18396 21364 18452 21534
rect 18396 21298 18452 21308
rect 18620 21252 18676 22094
rect 18732 21812 18788 22204
rect 18844 22194 18900 22204
rect 18956 22260 19012 22270
rect 18732 21746 18788 21756
rect 18956 21700 19012 22204
rect 18844 21644 19012 21700
rect 19180 21698 19236 23548
rect 19180 21646 19182 21698
rect 19234 21646 19236 21698
rect 18620 21186 18676 21196
rect 18732 21588 18788 21598
rect 17948 20916 18004 20926
rect 17836 20914 18004 20916
rect 17836 20862 17950 20914
rect 18002 20862 18004 20914
rect 17836 20860 18004 20862
rect 17948 20850 18004 20860
rect 18284 20916 18340 20926
rect 17388 20626 17444 20636
rect 17500 20804 17556 20814
rect 17052 20412 17332 20468
rect 15036 19406 15038 19458
rect 15090 19406 15092 19458
rect 15036 19394 15092 19406
rect 15708 19740 15988 19796
rect 14476 19294 14478 19346
rect 14530 19294 14532 19346
rect 14476 18452 14532 19294
rect 15148 19236 15204 19246
rect 15148 19142 15204 19180
rect 15036 19124 15092 19134
rect 15036 19030 15092 19068
rect 14588 18452 14644 18462
rect 15148 18452 15204 18462
rect 13916 18398 13918 18450
rect 13970 18398 13972 18450
rect 13916 18386 13972 18398
rect 14028 18450 15204 18452
rect 14028 18398 14590 18450
rect 14642 18398 15150 18450
rect 15202 18398 15204 18450
rect 14028 18396 15204 18398
rect 11788 18286 11790 18338
rect 11842 18286 11844 18338
rect 11788 18274 11844 18286
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 13468 16884 13524 16894
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16146 1988 16156
rect 13468 16210 13524 16828
rect 14028 16884 14084 18396
rect 14588 18386 14644 18396
rect 15148 18386 15204 18396
rect 15708 17666 15764 19740
rect 16268 18452 16324 18462
rect 15708 17614 15710 17666
rect 15762 17614 15764 17666
rect 15708 17602 15764 17614
rect 15820 17668 15876 17678
rect 15820 17574 15876 17612
rect 15932 17666 15988 17678
rect 15932 17614 15934 17666
rect 15986 17614 15988 17666
rect 14700 17444 14756 17454
rect 14700 16994 14756 17388
rect 15484 17444 15540 17454
rect 15484 17442 15652 17444
rect 15484 17390 15486 17442
rect 15538 17390 15652 17442
rect 15484 17388 15652 17390
rect 15484 17378 15540 17388
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 14028 16790 14084 16828
rect 13468 16158 13470 16210
rect 13522 16158 13524 16210
rect 13468 15428 13524 16158
rect 15596 16210 15652 17388
rect 15596 16158 15598 16210
rect 15650 16158 15652 16210
rect 15596 16146 15652 16158
rect 15708 15540 15764 15550
rect 15932 15540 15988 17614
rect 16268 17666 16324 18396
rect 16268 17614 16270 17666
rect 16322 17614 16324 17666
rect 16268 17602 16324 17614
rect 16716 17668 16772 17678
rect 16268 16884 16324 16894
rect 16268 16212 16324 16828
rect 16716 16884 16772 17612
rect 16828 17666 16884 20076
rect 17500 18450 17556 20748
rect 17500 18398 17502 18450
rect 17554 18398 17556 18450
rect 17500 18386 17556 18398
rect 17612 20580 17668 20590
rect 16828 17614 16830 17666
rect 16882 17614 16884 17666
rect 16828 17602 16884 17614
rect 17276 17666 17332 17678
rect 17276 17614 17278 17666
rect 17330 17614 17332 17666
rect 16940 17444 16996 17454
rect 16940 17350 16996 17388
rect 17276 16994 17332 17614
rect 17276 16942 17278 16994
rect 17330 16942 17332 16994
rect 17276 16930 17332 16942
rect 17500 16994 17556 17006
rect 17500 16942 17502 16994
rect 17554 16942 17556 16994
rect 16716 16818 16772 16828
rect 16828 16772 16884 16782
rect 17500 16772 17556 16942
rect 17612 16994 17668 20524
rect 17836 20578 17892 20590
rect 17836 20526 17838 20578
rect 17890 20526 17892 20578
rect 17724 18564 17780 18574
rect 17836 18564 17892 20526
rect 18060 20578 18116 20590
rect 18060 20526 18062 20578
rect 18114 20526 18116 20578
rect 18060 20244 18116 20526
rect 18284 20580 18340 20860
rect 18284 20486 18340 20524
rect 18060 20178 18116 20188
rect 18620 20244 18676 20254
rect 18732 20244 18788 21532
rect 18620 20242 18788 20244
rect 18620 20190 18622 20242
rect 18674 20190 18788 20242
rect 18620 20188 18788 20190
rect 18620 20178 18676 20188
rect 18844 19460 18900 21644
rect 19180 21634 19236 21646
rect 19292 23044 19348 23054
rect 19068 21588 19124 21598
rect 19068 20802 19124 21532
rect 19068 20750 19070 20802
rect 19122 20750 19124 20802
rect 19068 20738 19124 20750
rect 19180 21474 19236 21486
rect 19180 21422 19182 21474
rect 19234 21422 19236 21474
rect 18956 20692 19012 20702
rect 18956 20242 19012 20636
rect 18956 20190 18958 20242
rect 19010 20190 19012 20242
rect 18956 20178 19012 20190
rect 18844 19394 18900 19404
rect 19180 20020 19236 21422
rect 19292 20804 19348 22988
rect 19404 22260 19460 22270
rect 19404 21588 19460 22204
rect 19516 21812 19572 23884
rect 19628 23380 19684 24446
rect 20636 23940 20692 24670
rect 20972 24722 21028 24780
rect 20972 24670 20974 24722
rect 21026 24670 21028 24722
rect 20972 24658 21028 24670
rect 21196 24724 21252 25228
rect 21196 24630 21252 24668
rect 21980 24612 22036 24622
rect 21980 24610 22260 24612
rect 21980 24558 21982 24610
rect 22034 24558 22260 24610
rect 21980 24556 22260 24558
rect 21980 24546 22036 24556
rect 20636 23874 20692 23884
rect 21196 24276 21252 24286
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23314 19684 23324
rect 20188 23268 20244 23278
rect 19740 23044 19796 23054
rect 19740 22950 19796 22988
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21812 19684 21822
rect 20188 21812 20244 23212
rect 21084 23268 21140 23278
rect 21084 23174 21140 23212
rect 19516 21810 19684 21812
rect 19516 21758 19630 21810
rect 19682 21758 19684 21810
rect 19516 21756 19684 21758
rect 19628 21746 19684 21756
rect 20076 21756 20244 21812
rect 20412 23154 20468 23166
rect 20412 23102 20414 23154
rect 20466 23102 20468 23154
rect 19740 21700 19796 21710
rect 19740 21606 19796 21644
rect 19404 21532 19684 21588
rect 19404 21364 19460 21374
rect 19404 21026 19460 21308
rect 19404 20974 19406 21026
rect 19458 20974 19460 21026
rect 19404 20962 19460 20974
rect 19292 20748 19572 20804
rect 19292 20580 19348 20590
rect 19292 20486 19348 20524
rect 19404 20130 19460 20142
rect 19404 20078 19406 20130
rect 19458 20078 19460 20130
rect 19292 20020 19348 20030
rect 19180 20018 19348 20020
rect 19180 19966 19294 20018
rect 19346 19966 19348 20018
rect 19180 19964 19348 19966
rect 17724 18562 17892 18564
rect 17724 18510 17726 18562
rect 17778 18510 17892 18562
rect 17724 18508 17892 18510
rect 17724 18452 17780 18508
rect 17724 18386 17780 18396
rect 18732 18452 18788 18462
rect 18732 17106 18788 18396
rect 19180 18340 19236 19964
rect 19292 19954 19348 19964
rect 19180 18274 19236 18284
rect 19292 18562 19348 18574
rect 19292 18510 19294 18562
rect 19346 18510 19348 18562
rect 18732 17054 18734 17106
rect 18786 17054 18788 17106
rect 18732 17042 18788 17054
rect 18956 18116 19012 18126
rect 18956 17106 19012 18060
rect 19292 17332 19348 18510
rect 19404 18452 19460 20078
rect 19404 18386 19460 18396
rect 19516 18450 19572 20748
rect 19628 20130 19684 21532
rect 19964 21586 20020 21598
rect 19964 21534 19966 21586
rect 20018 21534 20020 21586
rect 19740 21252 19796 21262
rect 19740 20690 19796 21196
rect 19964 21140 20020 21534
rect 19964 21074 20020 21084
rect 19740 20638 19742 20690
rect 19794 20638 19796 20690
rect 19740 20626 19796 20638
rect 19964 20802 20020 20814
rect 19964 20750 19966 20802
rect 20018 20750 20020 20802
rect 19964 20692 20020 20750
rect 19964 20626 20020 20636
rect 20076 20580 20132 21756
rect 20188 21588 20244 21598
rect 20188 21494 20244 21532
rect 20412 21140 20468 23102
rect 20636 23156 20692 23166
rect 20636 21700 20692 23100
rect 21196 22596 21252 24220
rect 21756 23492 21812 23502
rect 21756 23378 21812 23436
rect 21756 23326 21758 23378
rect 21810 23326 21812 23378
rect 21308 23156 21364 23166
rect 21308 23062 21364 23100
rect 21644 23044 21700 23054
rect 21308 22596 21364 22606
rect 21196 22594 21364 22596
rect 21196 22542 21310 22594
rect 21362 22542 21364 22594
rect 21196 22540 21364 22542
rect 21308 22530 21364 22540
rect 21644 22594 21700 22988
rect 21644 22542 21646 22594
rect 21698 22542 21700 22594
rect 21644 22530 21700 22542
rect 21756 22484 21812 23326
rect 21868 23380 21924 23390
rect 21868 23286 21924 23324
rect 21980 23268 22036 23278
rect 21980 23174 22036 23212
rect 22204 22596 22260 24556
rect 22428 23268 22484 23278
rect 22428 23154 22484 23212
rect 22428 23102 22430 23154
rect 22482 23102 22484 23154
rect 22428 23090 22484 23102
rect 22540 23044 22596 25566
rect 23548 24724 23604 24734
rect 23548 24050 23604 24668
rect 24332 24724 24388 26126
rect 26236 26180 26292 26190
rect 26572 26180 26628 26238
rect 27916 26292 27972 26302
rect 26236 26178 26628 26180
rect 26236 26126 26238 26178
rect 26290 26126 26628 26178
rect 26236 26124 26628 26126
rect 27356 26178 27412 26190
rect 27356 26126 27358 26178
rect 27410 26126 27412 26178
rect 25340 25506 25396 25518
rect 25340 25454 25342 25506
rect 25394 25454 25396 25506
rect 24668 25394 24724 25406
rect 24668 25342 24670 25394
rect 24722 25342 24724 25394
rect 24668 24948 24724 25342
rect 24780 24948 24836 24958
rect 24668 24946 24836 24948
rect 24668 24894 24782 24946
rect 24834 24894 24836 24946
rect 24668 24892 24836 24894
rect 24780 24882 24836 24892
rect 24556 24834 24612 24846
rect 24556 24782 24558 24834
rect 24610 24782 24612 24834
rect 24332 24658 24388 24668
rect 24444 24722 24500 24734
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 23548 23998 23550 24050
rect 23602 23998 23604 24050
rect 23548 23986 23604 23998
rect 24108 24610 24164 24622
rect 24108 24558 24110 24610
rect 24162 24558 24164 24610
rect 22540 22978 22596 22988
rect 22652 23938 22708 23950
rect 22652 23886 22654 23938
rect 22706 23886 22708 23938
rect 22316 22596 22372 22606
rect 22204 22594 22372 22596
rect 22204 22542 22318 22594
rect 22370 22542 22372 22594
rect 22204 22540 22372 22542
rect 22316 22530 22372 22540
rect 21868 22484 21924 22494
rect 21756 22482 21924 22484
rect 21756 22430 21870 22482
rect 21922 22430 21924 22482
rect 21756 22428 21924 22430
rect 21868 22418 21924 22428
rect 22204 22260 22260 22270
rect 22204 22166 22260 22204
rect 22316 22148 22372 22158
rect 22316 22054 22372 22092
rect 21756 21812 21812 21822
rect 20636 21606 20692 21644
rect 21532 21698 21588 21710
rect 21532 21646 21534 21698
rect 21586 21646 21588 21698
rect 21532 21588 21588 21646
rect 20524 21364 20580 21374
rect 20524 21270 20580 21308
rect 20412 21084 20580 21140
rect 20412 20692 20468 20702
rect 20412 20598 20468 20636
rect 20524 20690 20580 21084
rect 21308 21028 21364 21038
rect 21308 20804 21364 20972
rect 20524 20638 20526 20690
rect 20578 20638 20580 20690
rect 20076 20524 20244 20580
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20244 20244 20524
rect 20076 20188 20244 20244
rect 19628 20078 19630 20130
rect 19682 20078 19684 20130
rect 19628 20066 19684 20078
rect 19964 20132 20020 20142
rect 19964 20038 20020 20076
rect 19852 20018 19908 20030
rect 19852 19966 19854 20018
rect 19906 19966 19908 20018
rect 19852 19572 19908 19966
rect 19964 19796 20020 19806
rect 19964 19702 20020 19740
rect 20076 19572 20132 20188
rect 20524 20132 20580 20638
rect 20524 20066 20580 20076
rect 21084 20802 21364 20804
rect 21084 20750 21310 20802
rect 21362 20750 21364 20802
rect 21084 20748 21364 20750
rect 21084 20130 21140 20748
rect 21308 20738 21364 20748
rect 21532 20188 21588 21532
rect 21756 21586 21812 21756
rect 21756 21534 21758 21586
rect 21810 21534 21812 21586
rect 21756 21522 21812 21534
rect 22204 21698 22260 21710
rect 22204 21646 22206 21698
rect 22258 21646 22260 21698
rect 22204 20804 22260 21646
rect 22428 21700 22484 21710
rect 22428 21586 22484 21644
rect 22428 21534 22430 21586
rect 22482 21534 22484 21586
rect 22428 21522 22484 21534
rect 22204 20356 22260 20748
rect 22204 20290 22260 20300
rect 22428 21140 22484 21150
rect 21084 20078 21086 20130
rect 21138 20078 21140 20130
rect 21084 20066 21140 20078
rect 21308 20132 21588 20188
rect 22316 20244 22372 20254
rect 19852 19516 20132 19572
rect 19852 19236 19908 19516
rect 19852 19170 19908 19180
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19516 18398 19518 18450
rect 19570 18398 19572 18450
rect 19516 18386 19572 18398
rect 19628 18340 19684 18350
rect 19516 17780 19572 17790
rect 19628 17780 19684 18284
rect 19740 18116 19796 18126
rect 19740 17890 19796 18060
rect 19740 17838 19742 17890
rect 19794 17838 19796 17890
rect 19740 17826 19796 17838
rect 19516 17778 19684 17780
rect 19516 17726 19518 17778
rect 19570 17726 19684 17778
rect 19516 17724 19684 17726
rect 19516 17714 19572 17724
rect 20076 17444 20132 17454
rect 20076 17442 20244 17444
rect 20076 17390 20078 17442
rect 20130 17390 20244 17442
rect 20076 17388 20244 17390
rect 20076 17378 20132 17388
rect 18956 17054 18958 17106
rect 19010 17054 19012 17106
rect 18956 17042 19012 17054
rect 19180 17276 19348 17332
rect 19836 17276 20100 17286
rect 17612 16942 17614 16994
rect 17666 16942 17668 16994
rect 17612 16930 17668 16942
rect 18284 16884 18340 16894
rect 16828 16770 17556 16772
rect 16828 16718 16830 16770
rect 16882 16718 17556 16770
rect 16828 16716 17556 16718
rect 17612 16772 17668 16782
rect 16268 16098 16324 16156
rect 16268 16046 16270 16098
rect 16322 16046 16324 16098
rect 16268 16034 16324 16046
rect 16604 16212 16660 16222
rect 15708 15538 15988 15540
rect 15708 15486 15710 15538
rect 15762 15486 15988 15538
rect 15708 15484 15988 15486
rect 15708 15474 15764 15484
rect 13468 15362 13524 15372
rect 15596 15428 15652 15438
rect 15596 15334 15652 15372
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 16604 14530 16660 16156
rect 16828 15148 16884 16716
rect 17052 16212 17108 16222
rect 17052 16118 17108 16156
rect 17500 16212 17556 16222
rect 17500 16118 17556 16156
rect 17612 15148 17668 16716
rect 18284 16658 18340 16828
rect 18508 16772 18564 16782
rect 18844 16772 18900 16782
rect 18508 16770 18676 16772
rect 18508 16718 18510 16770
rect 18562 16718 18676 16770
rect 18508 16716 18676 16718
rect 18508 16706 18564 16716
rect 18284 16606 18286 16658
rect 18338 16606 18340 16658
rect 18284 16100 18340 16606
rect 18620 16436 18676 16716
rect 18844 16678 18900 16716
rect 18620 16380 19124 16436
rect 18284 16034 18340 16044
rect 18956 16212 19012 16222
rect 16828 15092 17108 15148
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 16604 14466 16660 14478
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 16828 5236 16884 5246
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16828 800 16884 5180
rect 17052 5122 17108 15092
rect 17388 15092 17668 15148
rect 18956 15204 19012 16156
rect 19068 16210 19124 16380
rect 19068 16158 19070 16210
rect 19122 16158 19124 16210
rect 19068 16146 19124 16158
rect 19180 16100 19236 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 16882 20244 17388
rect 20188 16830 20190 16882
rect 20242 16830 20244 16882
rect 20188 16818 20244 16830
rect 20412 16994 20468 17006
rect 20412 16942 20414 16994
rect 20466 16942 20468 16994
rect 20412 16212 20468 16942
rect 21308 16322 21364 20132
rect 21980 20130 22036 20142
rect 21980 20078 21982 20130
rect 22034 20078 22036 20130
rect 21420 20018 21476 20030
rect 21420 19966 21422 20018
rect 21474 19966 21476 20018
rect 21420 19796 21476 19966
rect 21532 20020 21588 20030
rect 21532 19926 21588 19964
rect 21868 20018 21924 20030
rect 21868 19966 21870 20018
rect 21922 19966 21924 20018
rect 21868 19796 21924 19966
rect 21420 19740 21924 19796
rect 21308 16270 21310 16322
rect 21362 16270 21364 16322
rect 20412 16156 20692 16212
rect 19180 16034 19236 16044
rect 19852 16100 19908 16110
rect 19852 16006 19908 16044
rect 20188 16100 20244 16138
rect 20188 16034 20244 16044
rect 20636 16100 20692 16156
rect 20636 16098 21252 16100
rect 20636 16046 20638 16098
rect 20690 16046 21252 16098
rect 20636 16044 21252 16046
rect 20636 16034 20692 16044
rect 19292 15988 19348 15998
rect 19292 15894 19348 15932
rect 20412 15988 20468 15998
rect 20412 15894 20468 15932
rect 19068 15874 19124 15886
rect 19068 15822 19070 15874
rect 19122 15822 19124 15874
rect 19068 15652 19124 15822
rect 20188 15874 20244 15886
rect 20188 15822 20190 15874
rect 20242 15822 20244 15874
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19068 15596 19348 15652
rect 19836 15642 20100 15652
rect 17388 14642 17444 15092
rect 17388 14590 17390 14642
rect 17442 14590 17444 14642
rect 17388 14578 17444 14590
rect 18956 13746 19012 15148
rect 19292 15538 19348 15596
rect 20188 15540 20244 15822
rect 19292 15486 19294 15538
rect 19346 15486 19348 15538
rect 19292 15148 19348 15486
rect 19740 15484 20244 15540
rect 19628 15426 19684 15438
rect 19628 15374 19630 15426
rect 19682 15374 19684 15426
rect 19292 15092 19460 15148
rect 18956 13694 18958 13746
rect 19010 13694 19012 13746
rect 18956 13682 19012 13694
rect 19404 14644 19460 15092
rect 19516 14644 19572 14654
rect 19404 14642 19572 14644
rect 19404 14590 19518 14642
rect 19570 14590 19572 14642
rect 19404 14588 19572 14590
rect 18060 5236 18116 5246
rect 18060 5142 18116 5180
rect 17052 5070 17054 5122
rect 17106 5070 17108 5122
rect 17052 5058 17108 5070
rect 18844 3666 18900 3678
rect 18844 3614 18846 3666
rect 18898 3614 18900 3666
rect 18844 800 18900 3614
rect 19404 3556 19460 14588
rect 19516 14578 19572 14588
rect 19628 14420 19684 15374
rect 19516 14364 19684 14420
rect 19516 4340 19572 14364
rect 19740 14308 19796 15484
rect 21196 15428 21252 16044
rect 21308 15988 21364 16270
rect 21756 19234 21812 19246
rect 21756 19182 21758 19234
rect 21810 19182 21812 19234
rect 21420 16100 21476 16110
rect 21420 16006 21476 16044
rect 21308 15922 21364 15932
rect 21532 15874 21588 15886
rect 21532 15822 21534 15874
rect 21586 15822 21588 15874
rect 21308 15428 21364 15438
rect 21196 15426 21364 15428
rect 21196 15374 21310 15426
rect 21362 15374 21364 15426
rect 21196 15372 21364 15374
rect 21308 15362 21364 15372
rect 20524 15314 20580 15326
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 19964 15204 20020 15214
rect 19964 14642 20020 15148
rect 20524 15204 20580 15262
rect 20524 15138 20580 15148
rect 19964 14590 19966 14642
rect 20018 14590 20020 14642
rect 19964 14578 20020 14590
rect 19628 14252 19796 14308
rect 19628 13860 19684 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19740 13860 19796 13870
rect 19628 13858 19796 13860
rect 19628 13806 19742 13858
rect 19794 13806 19796 13858
rect 19628 13804 19796 13806
rect 19740 13794 19796 13804
rect 21532 13636 21588 15822
rect 21756 15204 21812 19182
rect 21868 18900 21924 19740
rect 21980 19348 22036 20078
rect 21980 19282 22036 19292
rect 22204 20018 22260 20030
rect 22204 19966 22206 20018
rect 22258 19966 22260 20018
rect 21868 18834 21924 18844
rect 22204 18452 22260 19966
rect 22316 19348 22372 20188
rect 22428 20242 22484 21084
rect 22428 20190 22430 20242
rect 22482 20190 22484 20242
rect 22428 20178 22484 20190
rect 22652 21140 22708 23886
rect 22764 23492 22820 23502
rect 22820 23436 22932 23492
rect 22764 23426 22820 23436
rect 22764 23266 22820 23278
rect 22764 23214 22766 23266
rect 22818 23214 22820 23266
rect 22764 23156 22820 23214
rect 22764 23090 22820 23100
rect 22764 21812 22820 21822
rect 22876 21812 22932 23436
rect 23100 23380 23156 23390
rect 23100 23286 23156 23324
rect 24108 23380 24164 24558
rect 24444 23492 24500 24670
rect 24444 23426 24500 23436
rect 24556 23828 24612 24782
rect 23660 23154 23716 23166
rect 23660 23102 23662 23154
rect 23714 23102 23716 23154
rect 23660 23044 23716 23102
rect 24108 23154 24164 23324
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 24108 23090 24164 23102
rect 24556 23268 24612 23772
rect 23660 22484 23716 22988
rect 22764 21810 22932 21812
rect 22764 21758 22766 21810
rect 22818 21758 22932 21810
rect 22764 21756 22932 21758
rect 23324 22428 23716 22484
rect 24220 23042 24276 23054
rect 24220 22990 24222 23042
rect 24274 22990 24276 23042
rect 22764 21746 22820 21756
rect 22428 19348 22484 19358
rect 22316 19346 22484 19348
rect 22316 19294 22430 19346
rect 22482 19294 22484 19346
rect 22316 19292 22484 19294
rect 22428 19282 22484 19292
rect 22204 18386 22260 18396
rect 22652 17666 22708 21084
rect 22988 21698 23044 21710
rect 22988 21646 22990 21698
rect 23042 21646 23044 21698
rect 22988 20916 23044 21646
rect 23100 21588 23156 21598
rect 23100 21586 23268 21588
rect 23100 21534 23102 21586
rect 23154 21534 23268 21586
rect 23100 21532 23268 21534
rect 23100 21522 23156 21532
rect 23100 20916 23156 20926
rect 22988 20860 23100 20916
rect 23100 20244 23156 20860
rect 22988 20242 23156 20244
rect 22988 20190 23102 20242
rect 23154 20190 23156 20242
rect 22988 20188 23156 20190
rect 22764 20020 22820 20030
rect 22764 18788 22820 19964
rect 22764 18722 22820 18732
rect 22876 19236 22932 19246
rect 22652 17614 22654 17666
rect 22706 17614 22708 17666
rect 22652 17602 22708 17614
rect 22764 18116 22820 18126
rect 22764 17106 22820 18060
rect 22764 17054 22766 17106
rect 22818 17054 22820 17106
rect 22764 17042 22820 17054
rect 22876 17108 22932 19180
rect 22988 18004 23044 20188
rect 23100 20178 23156 20188
rect 23100 18452 23156 18462
rect 23212 18452 23268 21532
rect 23324 20132 23380 22428
rect 24220 22372 24276 22990
rect 24556 22482 24612 23212
rect 24556 22430 24558 22482
rect 24610 22430 24612 22482
rect 24556 22418 24612 22430
rect 24892 24836 24948 24846
rect 24332 22372 24388 22382
rect 24220 22370 24500 22372
rect 24220 22318 24334 22370
rect 24386 22318 24500 22370
rect 24220 22316 24500 22318
rect 24332 22306 24388 22316
rect 23660 22260 23716 22270
rect 23660 22258 23940 22260
rect 23660 22206 23662 22258
rect 23714 22206 23940 22258
rect 23660 22204 23940 22206
rect 23660 22194 23716 22204
rect 23772 21698 23828 21710
rect 23772 21646 23774 21698
rect 23826 21646 23828 21698
rect 23436 21140 23492 21150
rect 23492 21084 23604 21140
rect 23436 21074 23492 21084
rect 23548 20914 23604 21084
rect 23548 20862 23550 20914
rect 23602 20862 23604 20914
rect 23548 20850 23604 20862
rect 23324 20018 23380 20076
rect 23324 19966 23326 20018
rect 23378 19966 23380 20018
rect 23324 19954 23380 19966
rect 23772 20020 23828 21646
rect 23884 20020 23940 22204
rect 24108 22258 24164 22270
rect 24108 22206 24110 22258
rect 24162 22206 24164 22258
rect 23996 21476 24052 21486
rect 24108 21476 24164 22206
rect 24444 21812 24500 22316
rect 24052 21420 24164 21476
rect 24220 21698 24276 21710
rect 24220 21646 24222 21698
rect 24274 21646 24276 21698
rect 23996 21410 24052 21420
rect 24220 20244 24276 21646
rect 24444 21586 24500 21756
rect 24668 21700 24724 21710
rect 24892 21700 24948 24780
rect 25340 24724 25396 25454
rect 25900 25284 25956 25294
rect 26236 25284 26292 26124
rect 27356 25730 27412 26126
rect 27356 25678 27358 25730
rect 27410 25678 27412 25730
rect 27356 25666 27412 25678
rect 27468 25508 27524 25518
rect 27468 25506 27860 25508
rect 27468 25454 27470 25506
rect 27522 25454 27860 25506
rect 27468 25452 27860 25454
rect 27468 25442 27524 25452
rect 26348 25284 26404 25294
rect 25900 25282 26740 25284
rect 25900 25230 25902 25282
rect 25954 25230 26350 25282
rect 26402 25230 26740 25282
rect 25900 25228 26740 25230
rect 25564 24724 25620 24734
rect 25900 24724 25956 25228
rect 26348 25218 26404 25228
rect 25396 24722 25956 24724
rect 25396 24670 25566 24722
rect 25618 24670 25956 24722
rect 25396 24668 25956 24670
rect 24668 21698 24948 21700
rect 24668 21646 24670 21698
rect 24722 21646 24948 21698
rect 24668 21644 24948 21646
rect 25228 21698 25284 21710
rect 25228 21646 25230 21698
rect 25282 21646 25284 21698
rect 24668 21634 24724 21644
rect 24444 21534 24446 21586
rect 24498 21534 24500 21586
rect 24444 21522 24500 21534
rect 25228 21476 25284 21646
rect 25228 21410 25284 21420
rect 24220 20178 24276 20188
rect 24332 20356 24388 20366
rect 24220 20020 24276 20030
rect 23884 20018 24276 20020
rect 23884 19966 24222 20018
rect 24274 19966 24276 20018
rect 23884 19964 24276 19966
rect 23772 19954 23828 19964
rect 23156 18396 23268 18452
rect 23436 18900 23492 18910
rect 23100 18386 23156 18396
rect 22988 17938 23044 17948
rect 23212 18228 23268 18238
rect 22988 17108 23044 17118
rect 22876 17106 23044 17108
rect 22876 17054 22990 17106
rect 23042 17054 23044 17106
rect 22876 17052 23044 17054
rect 22988 17042 23044 17052
rect 23212 17106 23268 18172
rect 23212 17054 23214 17106
rect 23266 17054 23268 17106
rect 23212 17042 23268 17054
rect 23324 17554 23380 17566
rect 23324 17502 23326 17554
rect 23378 17502 23380 17554
rect 22876 16772 22932 16782
rect 22876 16678 22932 16716
rect 23324 16098 23380 17502
rect 23324 16046 23326 16098
rect 23378 16046 23380 16098
rect 21756 15138 21812 15148
rect 22316 15204 22372 15214
rect 22316 13970 22372 15148
rect 23324 15204 23380 16046
rect 23324 15138 23380 15148
rect 23436 15202 23492 18844
rect 24108 18900 24164 18910
rect 24220 18900 24276 19964
rect 24164 18844 24276 18900
rect 24108 18834 24164 18844
rect 24332 18788 24388 20300
rect 24892 20244 24948 20254
rect 24444 20130 24500 20142
rect 24444 20078 24446 20130
rect 24498 20078 24500 20130
rect 24444 19460 24500 20078
rect 24444 19394 24500 19404
rect 24556 19348 24612 19358
rect 24556 19254 24612 19292
rect 24892 19236 24948 20188
rect 25340 20132 25396 24668
rect 25564 24658 25620 24668
rect 26348 24612 26404 24622
rect 26348 24518 26404 24556
rect 26684 23380 26740 25228
rect 27356 25282 27412 25294
rect 27692 25284 27748 25294
rect 27356 25230 27358 25282
rect 27410 25230 27412 25282
rect 27356 24836 27412 25230
rect 27356 24770 27412 24780
rect 27580 25282 27748 25284
rect 27580 25230 27694 25282
rect 27746 25230 27748 25282
rect 27580 25228 27748 25230
rect 27020 24612 27076 24622
rect 27020 24162 27076 24556
rect 27580 24388 27636 25228
rect 27692 25218 27748 25228
rect 27804 24500 27860 25452
rect 27916 25394 27972 26236
rect 37660 26292 37716 26302
rect 37660 26198 37716 26236
rect 29484 26178 29540 26190
rect 29484 26126 29486 26178
rect 29538 26126 29540 26178
rect 29260 25508 29316 25518
rect 29484 25508 29540 26126
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 39900 25620 39956 26126
rect 39900 25554 39956 25564
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 29260 25506 29540 25508
rect 29260 25454 29262 25506
rect 29314 25454 29540 25506
rect 29260 25452 29540 25454
rect 37660 25508 37716 25518
rect 27916 25342 27918 25394
rect 27970 25342 27972 25394
rect 27916 25172 27972 25342
rect 28028 25394 28084 25406
rect 28028 25342 28030 25394
rect 28082 25342 28084 25394
rect 28028 25284 28084 25342
rect 28028 25228 28644 25284
rect 27916 25116 28532 25172
rect 28364 24724 28420 24734
rect 27804 24444 28196 24500
rect 27020 24110 27022 24162
rect 27074 24110 27076 24162
rect 27020 24098 27076 24110
rect 27132 24332 27636 24388
rect 27132 23938 27188 24332
rect 27132 23886 27134 23938
rect 27186 23886 27188 23938
rect 27132 23874 27188 23886
rect 28140 23938 28196 24444
rect 28140 23886 28142 23938
rect 28194 23886 28196 23938
rect 28140 23874 28196 23886
rect 27020 23828 27076 23838
rect 27020 23734 27076 23772
rect 28364 23826 28420 24668
rect 28476 24610 28532 25116
rect 28476 24558 28478 24610
rect 28530 24558 28532 24610
rect 28476 24546 28532 24558
rect 28476 23940 28532 23950
rect 28588 23940 28644 25228
rect 29260 24724 29316 25452
rect 37660 25414 37716 25452
rect 29484 25284 29540 25294
rect 29484 25190 29540 25228
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 29260 24658 29316 24668
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 28476 23938 28588 23940
rect 28476 23886 28478 23938
rect 28530 23886 28588 23938
rect 28476 23884 28588 23886
rect 28476 23874 28532 23884
rect 28588 23846 28644 23884
rect 28924 23940 28980 23950
rect 28364 23774 28366 23826
rect 28418 23774 28420 23826
rect 28364 23762 28420 23774
rect 28028 23716 28084 23726
rect 26796 23380 26852 23390
rect 26684 23378 27188 23380
rect 26684 23326 26798 23378
rect 26850 23326 27188 23378
rect 26684 23324 27188 23326
rect 26796 23286 26852 23324
rect 27132 23154 27188 23324
rect 27132 23102 27134 23154
rect 27186 23102 27188 23154
rect 27132 23090 27188 23102
rect 27916 23042 27972 23054
rect 27916 22990 27918 23042
rect 27970 22990 27972 23042
rect 27916 22594 27972 22990
rect 27916 22542 27918 22594
rect 27970 22542 27972 22594
rect 27916 22530 27972 22542
rect 28028 22370 28084 23660
rect 28028 22318 28030 22370
rect 28082 22318 28084 22370
rect 28028 22306 28084 22318
rect 27916 22148 27972 22158
rect 27916 22054 27972 22092
rect 27804 21698 27860 21710
rect 27804 21646 27806 21698
rect 27858 21646 27860 21698
rect 25564 21588 25620 21598
rect 25564 21586 25844 21588
rect 25564 21534 25566 21586
rect 25618 21534 25844 21586
rect 25564 21532 25844 21534
rect 25564 21522 25620 21532
rect 25340 20130 25732 20132
rect 25340 20078 25342 20130
rect 25394 20078 25732 20130
rect 25340 20076 25732 20078
rect 25340 20066 25396 20076
rect 25676 20018 25732 20076
rect 25676 19966 25678 20018
rect 25730 19966 25732 20018
rect 25676 19954 25732 19966
rect 25676 19348 25732 19358
rect 25788 19348 25844 21532
rect 27580 21586 27636 21598
rect 27580 21534 27582 21586
rect 27634 21534 27636 21586
rect 27580 20188 27636 21534
rect 27804 21588 27860 21646
rect 27804 21522 27860 21532
rect 27916 21586 27972 21598
rect 27916 21534 27918 21586
rect 27970 21534 27972 21586
rect 27916 20468 27972 21534
rect 27916 20402 27972 20412
rect 28588 21588 28644 21598
rect 26908 20132 27636 20188
rect 26460 19908 26516 19918
rect 26460 19906 26628 19908
rect 26460 19854 26462 19906
rect 26514 19854 26628 19906
rect 26460 19852 26628 19854
rect 26460 19842 26516 19852
rect 26124 19796 26180 19806
rect 26124 19458 26180 19740
rect 26124 19406 26126 19458
rect 26178 19406 26180 19458
rect 26124 19394 26180 19406
rect 26348 19460 26404 19470
rect 26348 19366 26404 19404
rect 25732 19292 25844 19348
rect 26572 19346 26628 19852
rect 26908 19458 26964 20132
rect 28588 19906 28644 21532
rect 28588 19854 28590 19906
rect 28642 19854 28644 19906
rect 28588 19842 28644 19854
rect 28812 20468 28868 20478
rect 28812 19908 28868 20412
rect 28924 20188 28980 23884
rect 29372 23940 29428 23950
rect 29372 23846 29428 23884
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 29036 23716 29092 23726
rect 29036 23622 29092 23660
rect 29260 23716 29316 23726
rect 29260 23622 29316 23660
rect 30044 23716 30100 23726
rect 30044 23042 30100 23660
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 30044 22990 30046 23042
rect 30098 22990 30100 23042
rect 30044 22978 30100 22990
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21362 40068 21374
rect 40012 21310 40014 21362
rect 40066 21310 40068 21362
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 40012 20916 40068 21310
rect 40012 20850 40068 20860
rect 30044 20468 30100 20478
rect 28924 20132 29652 20188
rect 28924 20130 28980 20132
rect 28924 20078 28926 20130
rect 28978 20078 28980 20130
rect 28924 20066 28980 20078
rect 29596 20130 29652 20132
rect 29596 20078 29598 20130
rect 29650 20078 29652 20130
rect 29596 20066 29652 20078
rect 29708 20132 29764 20142
rect 29764 20076 29876 20132
rect 29708 20038 29764 20076
rect 29148 20018 29204 20030
rect 29148 19966 29150 20018
rect 29202 19966 29204 20018
rect 29148 19908 29204 19966
rect 28812 19852 29204 19908
rect 29708 19794 29764 19806
rect 29708 19742 29710 19794
rect 29762 19742 29764 19794
rect 26908 19406 26910 19458
rect 26962 19406 26964 19458
rect 26908 19394 26964 19406
rect 27244 19572 27300 19582
rect 26572 19294 26574 19346
rect 26626 19294 26628 19346
rect 25676 19254 25732 19292
rect 26572 19282 26628 19294
rect 24892 19122 24948 19180
rect 26684 19236 26740 19246
rect 26684 19142 26740 19180
rect 27244 19234 27300 19516
rect 29372 19572 29428 19582
rect 27244 19182 27246 19234
rect 27298 19182 27300 19234
rect 27244 19170 27300 19182
rect 27804 19236 27860 19246
rect 27804 19142 27860 19180
rect 29372 19234 29428 19516
rect 29372 19182 29374 19234
rect 29426 19182 29428 19234
rect 29372 19170 29428 19182
rect 29708 19234 29764 19742
rect 29708 19182 29710 19234
rect 29762 19182 29764 19234
rect 29708 19170 29764 19182
rect 24892 19070 24894 19122
rect 24946 19070 24948 19122
rect 24892 19058 24948 19070
rect 25228 19012 25284 19022
rect 25564 19012 25620 19022
rect 25228 19010 25620 19012
rect 25228 18958 25230 19010
rect 25282 18958 25566 19010
rect 25618 18958 25620 19010
rect 25228 18956 25620 18958
rect 25228 18946 25284 18956
rect 24220 18732 24388 18788
rect 25228 18788 25284 18798
rect 23884 18562 23940 18574
rect 23884 18510 23886 18562
rect 23938 18510 23940 18562
rect 23548 18452 23604 18462
rect 23548 18358 23604 18396
rect 23884 18452 23940 18510
rect 24220 18562 24276 18732
rect 24220 18510 24222 18562
rect 24274 18510 24276 18562
rect 24220 18498 24276 18510
rect 24332 18564 24388 18574
rect 24332 18470 24388 18508
rect 25116 18564 25172 18574
rect 23884 18386 23940 18396
rect 24332 18228 24388 18238
rect 25116 18228 25172 18508
rect 25228 18562 25284 18732
rect 25340 18674 25396 18956
rect 25564 18946 25620 18956
rect 26460 19012 26516 19022
rect 25340 18622 25342 18674
rect 25394 18622 25396 18674
rect 25340 18610 25396 18622
rect 25228 18510 25230 18562
rect 25282 18510 25284 18562
rect 25228 18498 25284 18510
rect 25900 18340 25956 18350
rect 25788 18284 25900 18340
rect 25340 18228 25396 18238
rect 25116 18172 25284 18228
rect 24332 18134 24388 18172
rect 23660 18004 23716 18014
rect 23660 16882 23716 17948
rect 23660 16830 23662 16882
rect 23714 16830 23716 16882
rect 23660 16818 23716 16830
rect 24556 16884 24612 16894
rect 23884 16772 23940 16782
rect 23884 16678 23940 16716
rect 24220 16660 24276 16670
rect 23996 16658 24276 16660
rect 23996 16606 24222 16658
rect 24274 16606 24276 16658
rect 23996 16604 24276 16606
rect 23884 15316 23940 15326
rect 23996 15316 24052 16604
rect 24220 16594 24276 16604
rect 24108 15986 24164 15998
rect 24108 15934 24110 15986
rect 24162 15934 24164 15986
rect 24108 15538 24164 15934
rect 24108 15486 24110 15538
rect 24162 15486 24164 15538
rect 24108 15474 24164 15486
rect 23884 15314 24052 15316
rect 23884 15262 23886 15314
rect 23938 15262 24052 15314
rect 23884 15260 24052 15262
rect 23884 15250 23940 15260
rect 23436 15150 23438 15202
rect 23490 15150 23492 15202
rect 23436 15138 23492 15150
rect 24556 15204 24612 16828
rect 25228 15540 25284 18172
rect 25340 18134 25396 18172
rect 25340 16884 25396 16894
rect 25340 16790 25396 16828
rect 25788 16884 25844 18284
rect 25900 18246 25956 18284
rect 26460 16994 26516 18956
rect 27356 19012 27412 19022
rect 27356 18918 27412 18956
rect 27468 19010 27524 19022
rect 27468 18958 27470 19010
rect 27522 18958 27524 19010
rect 27020 18450 27076 18462
rect 27020 18398 27022 18450
rect 27074 18398 27076 18450
rect 26572 18340 26628 18350
rect 26572 18246 26628 18284
rect 27020 18340 27076 18398
rect 27468 18452 27524 18958
rect 29148 19010 29204 19022
rect 29148 18958 29150 19010
rect 29202 18958 29204 19010
rect 27468 18386 27524 18396
rect 27692 18564 27748 18574
rect 27692 18450 27748 18508
rect 27692 18398 27694 18450
rect 27746 18398 27748 18450
rect 27692 18386 27748 18398
rect 27020 18274 27076 18284
rect 29148 18228 29204 18958
rect 29260 19010 29316 19022
rect 29260 18958 29262 19010
rect 29314 18958 29316 19010
rect 29260 18564 29316 18958
rect 29260 18498 29316 18508
rect 29820 18338 29876 20076
rect 30044 19234 30100 20412
rect 37660 20132 37716 20142
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 30044 19182 30046 19234
rect 30098 19182 30100 19234
rect 30044 19170 30100 19182
rect 30380 19236 30436 19246
rect 30380 19142 30436 19180
rect 37660 19234 37716 20076
rect 37660 19182 37662 19234
rect 37714 19182 37716 19234
rect 37660 19170 37716 19182
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 29820 18286 29822 18338
rect 29874 18286 29876 18338
rect 29820 18274 29876 18286
rect 30156 19010 30212 19022
rect 30156 18958 30158 19010
rect 30210 18958 30212 19010
rect 30156 18452 30212 18958
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 29148 18162 29204 18172
rect 26460 16942 26462 16994
rect 26514 16942 26516 16994
rect 26460 16930 26516 16942
rect 28588 18116 28644 18126
rect 25788 16790 25844 16828
rect 26908 16884 26964 16894
rect 26908 16210 26964 16828
rect 28588 16770 28644 18060
rect 30156 18116 30212 18396
rect 37660 18452 37716 18462
rect 37660 18358 37716 18396
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 30156 18050 30212 18060
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 28588 16718 28590 16770
rect 28642 16718 28644 16770
rect 28588 16706 28644 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 26908 16158 26910 16210
rect 26962 16158 26964 16210
rect 26908 16146 26964 16158
rect 26348 15874 26404 15886
rect 26348 15822 26350 15874
rect 26402 15822 26404 15874
rect 25228 15446 25284 15484
rect 25900 15540 25956 15550
rect 25900 15446 25956 15484
rect 26348 15540 26404 15822
rect 26348 15474 26404 15484
rect 24556 15138 24612 15148
rect 25564 15426 25620 15438
rect 25564 15374 25566 15426
rect 25618 15374 25620 15426
rect 25564 15148 25620 15374
rect 26236 15428 26292 15438
rect 26236 15334 26292 15372
rect 28588 15428 28644 15438
rect 27020 15316 27076 15326
rect 25564 15092 25844 15148
rect 22316 13918 22318 13970
rect 22370 13918 22372 13970
rect 22316 13906 22372 13918
rect 21868 13636 21924 13646
rect 21532 13634 21924 13636
rect 21532 13582 21870 13634
rect 21922 13582 21924 13634
rect 21532 13580 21924 13582
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19740 4340 19796 4350
rect 19516 4338 19796 4340
rect 19516 4286 19742 4338
rect 19794 4286 19796 4338
rect 19516 4284 19796 4286
rect 19740 4274 19796 4284
rect 19964 4116 20020 4126
rect 19740 3556 19796 3566
rect 19404 3554 19796 3556
rect 19404 3502 19742 3554
rect 19794 3502 19796 3554
rect 19404 3500 19796 3502
rect 19740 3490 19796 3500
rect 19964 3388 20020 4060
rect 20748 4116 20804 4126
rect 20748 4022 20804 4060
rect 19516 3332 20020 3388
rect 21532 3668 21588 3678
rect 19516 800 19572 3332
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 21532 800 21588 3612
rect 21756 3554 21812 13580
rect 21868 13570 21924 13580
rect 25788 4338 25844 15092
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 25564 4116 25620 4126
rect 22428 3668 22484 3678
rect 22428 3574 22484 3612
rect 24780 3666 24836 3678
rect 24780 3614 24782 3666
rect 24834 3614 24836 3666
rect 21756 3502 21758 3554
rect 21810 3502 21812 3554
rect 21756 3490 21812 3502
rect 24780 3388 24836 3614
rect 24220 3332 24836 3388
rect 24220 800 24276 3332
rect 25564 800 25620 4060
rect 26796 4116 26852 4126
rect 26796 4022 26852 4060
rect 26236 3668 26292 3678
rect 26236 800 26292 3612
rect 27020 3554 27076 15260
rect 27020 3502 27022 3554
rect 27074 3502 27076 3554
rect 27020 3490 27076 3502
rect 28588 3554 28644 15372
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 16800 0 16912 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 21504 0 21616 800
rect 24192 0 24304 800
rect 25536 0 25648 800
rect 26208 0 26320 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 16156 37884 16212 37940
rect 16940 37938 16996 37940
rect 16940 37886 16942 37938
rect 16942 37886 16994 37938
rect 16994 37886 16996 37938
rect 16940 37884 16996 37886
rect 17500 37436 17556 37492
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4172 26236 4228 26292
rect 1932 24892 1988 24948
rect 1932 23548 1988 23604
rect 1932 22482 1988 22484
rect 1932 22430 1934 22482
rect 1934 22430 1986 22482
rect 1986 22430 1988 22482
rect 1932 22428 1988 22430
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 11788 25452 11844 25508
rect 11788 24892 11844 24948
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 12684 24220 12740 24276
rect 4284 22988 4340 23044
rect 11564 23100 11620 23156
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4284 22370 4340 22372
rect 4284 22318 4286 22370
rect 4286 22318 4338 22370
rect 4338 22318 4340 22370
rect 4284 22316 4340 22318
rect 11004 22316 11060 22372
rect 13916 25228 13972 25284
rect 14700 25228 14756 25284
rect 13804 25116 13860 25172
rect 16604 25618 16660 25620
rect 16604 25566 16606 25618
rect 16606 25566 16658 25618
rect 16658 25566 16660 25618
rect 16604 25564 16660 25566
rect 14812 25004 14868 25060
rect 15372 25116 15428 25172
rect 15260 24946 15316 24948
rect 15260 24894 15262 24946
rect 15262 24894 15314 24946
rect 15314 24894 15316 24946
rect 15260 24892 15316 24894
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18508 37490 18564 37492
rect 18508 37438 18510 37490
rect 18510 37438 18562 37490
rect 18562 37438 18564 37490
rect 18508 37436 18564 37438
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 20860 38220 20916 38276
rect 22092 38274 22148 38276
rect 22092 38222 22094 38274
rect 22094 38222 22146 38274
rect 22146 38222 22148 38274
rect 22092 38220 22148 38222
rect 20188 37436 20244 37492
rect 20860 37266 20916 37268
rect 20860 37214 20862 37266
rect 20862 37214 20914 37266
rect 20914 37214 20916 37266
rect 20860 37212 20916 37214
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17612 25564 17668 25620
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 18844 25564 18900 25620
rect 17948 25228 18004 25284
rect 17724 25004 17780 25060
rect 13468 24220 13524 24276
rect 13804 23938 13860 23940
rect 13804 23886 13806 23938
rect 13806 23886 13858 23938
rect 13858 23886 13860 23938
rect 13804 23884 13860 23886
rect 15036 24722 15092 24724
rect 15036 24670 15038 24722
rect 15038 24670 15090 24722
rect 15090 24670 15092 24722
rect 15036 24668 15092 24670
rect 14924 23884 14980 23940
rect 14028 23548 14084 23604
rect 14812 23324 14868 23380
rect 14924 23436 14980 23492
rect 17500 24722 17556 24724
rect 17500 24670 17502 24722
rect 17502 24670 17554 24722
rect 17554 24670 17556 24722
rect 17500 24668 17556 24670
rect 15708 23660 15764 23716
rect 17388 23660 17444 23716
rect 15932 23378 15988 23380
rect 15932 23326 15934 23378
rect 15934 23326 15986 23378
rect 15986 23326 15988 23378
rect 15932 23324 15988 23326
rect 15036 23154 15092 23156
rect 15036 23102 15038 23154
rect 15038 23102 15090 23154
rect 15090 23102 15092 23154
rect 15036 23100 15092 23102
rect 14252 22370 14308 22372
rect 14252 22318 14254 22370
rect 14254 22318 14306 22370
rect 14306 22318 14308 22370
rect 14252 22316 14308 22318
rect 12908 22258 12964 22260
rect 12908 22206 12910 22258
rect 12910 22206 12962 22258
rect 12962 22206 12964 22258
rect 12908 22204 12964 22206
rect 14140 22258 14196 22260
rect 14140 22206 14142 22258
rect 14142 22206 14194 22258
rect 14194 22206 14196 22258
rect 14140 22204 14196 22206
rect 15260 23154 15316 23156
rect 15260 23102 15262 23154
rect 15262 23102 15314 23154
rect 15314 23102 15316 23154
rect 15260 23100 15316 23102
rect 16604 23100 16660 23156
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 14588 21084 14644 21140
rect 4172 20972 4228 21028
rect 1932 20188 1988 20244
rect 13804 20636 13860 20692
rect 11788 20076 11844 20132
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 11340 19964 11396 20020
rect 4172 19852 4228 19908
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 11788 19068 11844 19124
rect 16604 22316 16660 22372
rect 15484 22204 15540 22260
rect 15260 20802 15316 20804
rect 15260 20750 15262 20802
rect 15262 20750 15314 20802
rect 15314 20750 15316 20802
rect 15260 20748 15316 20750
rect 14924 20636 14980 20692
rect 16156 22204 16212 22260
rect 15932 21084 15988 21140
rect 14588 20242 14644 20244
rect 14588 20190 14590 20242
rect 14590 20190 14642 20242
rect 14642 20190 14644 20242
rect 14588 20188 14644 20190
rect 15260 20076 15316 20132
rect 13916 19852 13972 19908
rect 14812 20018 14868 20020
rect 14812 19966 14814 20018
rect 14814 19966 14866 20018
rect 14866 19966 14868 20018
rect 14812 19964 14868 19966
rect 15036 19964 15092 20020
rect 15708 20018 15764 20020
rect 15708 19966 15710 20018
rect 15710 19966 15762 20018
rect 15762 19966 15764 20018
rect 15708 19964 15764 19966
rect 15596 19906 15652 19908
rect 15596 19854 15598 19906
rect 15598 19854 15650 19906
rect 15650 19854 15652 19906
rect 15596 19852 15652 19854
rect 16940 22258 16996 22260
rect 16940 22206 16942 22258
rect 16942 22206 16994 22258
rect 16994 22206 16996 22258
rect 16940 22204 16996 22206
rect 17276 21644 17332 21700
rect 17164 21532 17220 21588
rect 16492 20860 16548 20916
rect 16716 21084 16772 21140
rect 16716 20802 16772 20804
rect 16716 20750 16718 20802
rect 16718 20750 16770 20802
rect 16770 20750 16772 20802
rect 16716 20748 16772 20750
rect 16044 20188 16100 20244
rect 17836 24722 17892 24724
rect 17836 24670 17838 24722
rect 17838 24670 17890 24722
rect 17890 24670 17892 24722
rect 17836 24668 17892 24670
rect 17500 23548 17556 23604
rect 17612 22370 17668 22372
rect 17612 22318 17614 22370
rect 17614 22318 17666 22370
rect 17666 22318 17668 22370
rect 17612 22316 17668 22318
rect 17836 22370 17892 22372
rect 17836 22318 17838 22370
rect 17838 22318 17890 22370
rect 17890 22318 17892 22370
rect 17836 22316 17892 22318
rect 21644 37212 21700 37268
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 40236 36370 40292 36372
rect 40236 36318 40238 36370
rect 40238 36318 40290 36370
rect 40290 36318 40292 36370
rect 40236 36316 40292 36318
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19404 25228 19460 25284
rect 19964 25282 20020 25284
rect 19964 25230 19966 25282
rect 19966 25230 20018 25282
rect 20018 25230 20020 25282
rect 19964 25228 20020 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20972 25228 21028 25284
rect 18956 24834 19012 24836
rect 18956 24782 18958 24834
rect 18958 24782 19010 24834
rect 19010 24782 19012 24834
rect 18956 24780 19012 24782
rect 20972 24780 21028 24836
rect 18732 24668 18788 24724
rect 18060 22258 18116 22260
rect 18060 22206 18062 22258
rect 18062 22206 18114 22258
rect 18114 22206 18116 22258
rect 18060 22204 18116 22206
rect 18732 23660 18788 23716
rect 19180 23938 19236 23940
rect 19180 23886 19182 23938
rect 19182 23886 19234 23938
rect 19234 23886 19236 23938
rect 19180 23884 19236 23886
rect 19740 24722 19796 24724
rect 19740 24670 19742 24722
rect 19742 24670 19794 24722
rect 19794 24670 19796 24722
rect 19740 24668 19796 24670
rect 19516 24220 19572 24276
rect 19516 23884 19572 23940
rect 18956 22988 19012 23044
rect 19180 23548 19236 23604
rect 18396 22258 18452 22260
rect 18396 22206 18398 22258
rect 18398 22206 18450 22258
rect 18450 22206 18452 22258
rect 18396 22204 18452 22206
rect 18172 22146 18228 22148
rect 18172 22094 18174 22146
rect 18174 22094 18226 22146
rect 18226 22094 18228 22146
rect 18172 22092 18228 22094
rect 17724 21810 17780 21812
rect 17724 21758 17726 21810
rect 17726 21758 17778 21810
rect 17778 21758 17780 21810
rect 17724 21756 17780 21758
rect 18396 21756 18452 21812
rect 18396 21308 18452 21364
rect 18956 22204 19012 22260
rect 18732 21756 18788 21812
rect 18620 21196 18676 21252
rect 18732 21586 18788 21588
rect 18732 21534 18734 21586
rect 18734 21534 18786 21586
rect 18786 21534 18788 21586
rect 18732 21532 18788 21534
rect 18284 20860 18340 20916
rect 17388 20636 17444 20692
rect 17500 20748 17556 20804
rect 16828 20076 16884 20132
rect 15148 19234 15204 19236
rect 15148 19182 15150 19234
rect 15150 19182 15202 19234
rect 15202 19182 15204 19234
rect 15148 19180 15204 19182
rect 15036 19122 15092 19124
rect 15036 19070 15038 19122
rect 15038 19070 15090 19122
rect 15090 19070 15092 19122
rect 15036 19068 15092 19070
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 13468 16828 13524 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 16156 1988 16212
rect 16268 18396 16324 18452
rect 15820 17666 15876 17668
rect 15820 17614 15822 17666
rect 15822 17614 15874 17666
rect 15874 17614 15876 17666
rect 15820 17612 15876 17614
rect 14700 17388 14756 17444
rect 14028 16882 14084 16884
rect 14028 16830 14030 16882
rect 14030 16830 14082 16882
rect 14082 16830 14084 16882
rect 14028 16828 14084 16830
rect 16716 17666 16772 17668
rect 16716 17614 16718 17666
rect 16718 17614 16770 17666
rect 16770 17614 16772 17666
rect 16716 17612 16772 17614
rect 16268 16828 16324 16884
rect 17612 20524 17668 20580
rect 16940 17442 16996 17444
rect 16940 17390 16942 17442
rect 16942 17390 16994 17442
rect 16994 17390 16996 17442
rect 16940 17388 16996 17390
rect 16716 16828 16772 16884
rect 18284 20578 18340 20580
rect 18284 20526 18286 20578
rect 18286 20526 18338 20578
rect 18338 20526 18340 20578
rect 18284 20524 18340 20526
rect 18060 20188 18116 20244
rect 19292 22988 19348 23044
rect 19068 21532 19124 21588
rect 18956 20636 19012 20692
rect 18844 19404 18900 19460
rect 19404 22204 19460 22260
rect 21196 24722 21252 24724
rect 21196 24670 21198 24722
rect 21198 24670 21250 24722
rect 21250 24670 21252 24722
rect 21196 24668 21252 24670
rect 20636 23884 20692 23940
rect 21196 24220 21252 24276
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19628 23324 19684 23380
rect 20188 23212 20244 23268
rect 19740 23042 19796 23044
rect 19740 22990 19742 23042
rect 19742 22990 19794 23042
rect 19794 22990 19796 23042
rect 19740 22988 19796 22990
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21084 23266 21140 23268
rect 21084 23214 21086 23266
rect 21086 23214 21138 23266
rect 21138 23214 21140 23266
rect 21084 23212 21140 23214
rect 19740 21698 19796 21700
rect 19740 21646 19742 21698
rect 19742 21646 19794 21698
rect 19794 21646 19796 21698
rect 19740 21644 19796 21646
rect 19404 21308 19460 21364
rect 19292 20578 19348 20580
rect 19292 20526 19294 20578
rect 19294 20526 19346 20578
rect 19346 20526 19348 20578
rect 19292 20524 19348 20526
rect 17724 18396 17780 18452
rect 18732 18396 18788 18452
rect 19180 18284 19236 18340
rect 18956 18060 19012 18116
rect 19404 18396 19460 18452
rect 19740 21196 19796 21252
rect 19964 21084 20020 21140
rect 19964 20636 20020 20692
rect 20188 21586 20244 21588
rect 20188 21534 20190 21586
rect 20190 21534 20242 21586
rect 20242 21534 20244 21586
rect 20188 21532 20244 21534
rect 20636 23154 20692 23156
rect 20636 23102 20638 23154
rect 20638 23102 20690 23154
rect 20690 23102 20692 23154
rect 20636 23100 20692 23102
rect 21756 23436 21812 23492
rect 21308 23154 21364 23156
rect 21308 23102 21310 23154
rect 21310 23102 21362 23154
rect 21362 23102 21364 23154
rect 21308 23100 21364 23102
rect 21644 22988 21700 23044
rect 21868 23378 21924 23380
rect 21868 23326 21870 23378
rect 21870 23326 21922 23378
rect 21922 23326 21924 23378
rect 21868 23324 21924 23326
rect 21980 23266 22036 23268
rect 21980 23214 21982 23266
rect 21982 23214 22034 23266
rect 22034 23214 22036 23266
rect 21980 23212 22036 23214
rect 22428 23212 22484 23268
rect 23548 24668 23604 24724
rect 27916 26236 27972 26292
rect 24332 24668 24388 24724
rect 22540 22988 22596 23044
rect 22204 22258 22260 22260
rect 22204 22206 22206 22258
rect 22206 22206 22258 22258
rect 22258 22206 22260 22258
rect 22204 22204 22260 22206
rect 22316 22146 22372 22148
rect 22316 22094 22318 22146
rect 22318 22094 22370 22146
rect 22370 22094 22372 22146
rect 22316 22092 22372 22094
rect 21756 21756 21812 21812
rect 20636 21698 20692 21700
rect 20636 21646 20638 21698
rect 20638 21646 20690 21698
rect 20690 21646 20692 21698
rect 20636 21644 20692 21646
rect 21532 21532 21588 21588
rect 20524 21362 20580 21364
rect 20524 21310 20526 21362
rect 20526 21310 20578 21362
rect 20578 21310 20580 21362
rect 20524 21308 20580 21310
rect 20412 20690 20468 20692
rect 20412 20638 20414 20690
rect 20414 20638 20466 20690
rect 20466 20638 20468 20690
rect 20412 20636 20468 20638
rect 21308 20972 21364 21028
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19964 20130 20020 20132
rect 19964 20078 19966 20130
rect 19966 20078 20018 20130
rect 20018 20078 20020 20130
rect 19964 20076 20020 20078
rect 19964 19794 20020 19796
rect 19964 19742 19966 19794
rect 19966 19742 20018 19794
rect 20018 19742 20020 19794
rect 19964 19740 20020 19742
rect 20524 20076 20580 20132
rect 22428 21644 22484 21700
rect 22204 20748 22260 20804
rect 22204 20300 22260 20356
rect 22428 21084 22484 21140
rect 22316 20188 22372 20244
rect 19852 19180 19908 19236
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18284 19684 18340
rect 19740 18060 19796 18116
rect 18284 16828 18340 16884
rect 17612 16716 17668 16772
rect 16268 16156 16324 16212
rect 16604 16156 16660 16212
rect 13468 15372 13524 15428
rect 15596 15426 15652 15428
rect 15596 15374 15598 15426
rect 15598 15374 15650 15426
rect 15650 15374 15652 15426
rect 15596 15372 15652 15374
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 17052 16210 17108 16212
rect 17052 16158 17054 16210
rect 17054 16158 17106 16210
rect 17106 16158 17108 16210
rect 17052 16156 17108 16158
rect 17500 16210 17556 16212
rect 17500 16158 17502 16210
rect 17502 16158 17554 16210
rect 17554 16158 17556 16210
rect 17500 16156 17556 16158
rect 18844 16770 18900 16772
rect 18844 16718 18846 16770
rect 18846 16718 18898 16770
rect 18898 16718 18900 16770
rect 18844 16716 18900 16718
rect 18284 16044 18340 16100
rect 18956 16156 19012 16212
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 16828 5180 16884 5236
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 21532 20018 21588 20020
rect 21532 19966 21534 20018
rect 21534 19966 21586 20018
rect 21586 19966 21588 20018
rect 21532 19964 21588 19966
rect 19180 16044 19236 16100
rect 19852 16098 19908 16100
rect 19852 16046 19854 16098
rect 19854 16046 19906 16098
rect 19906 16046 19908 16098
rect 19852 16044 19908 16046
rect 20188 16098 20244 16100
rect 20188 16046 20190 16098
rect 20190 16046 20242 16098
rect 20242 16046 20244 16098
rect 20188 16044 20244 16046
rect 19292 15986 19348 15988
rect 19292 15934 19294 15986
rect 19294 15934 19346 15986
rect 19346 15934 19348 15986
rect 19292 15932 19348 15934
rect 20412 15986 20468 15988
rect 20412 15934 20414 15986
rect 20414 15934 20466 15986
rect 20466 15934 20468 15986
rect 20412 15932 20468 15934
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18956 15148 19012 15204
rect 18060 5234 18116 5236
rect 18060 5182 18062 5234
rect 18062 5182 18114 5234
rect 18114 5182 18116 5234
rect 18060 5180 18116 5182
rect 21420 16098 21476 16100
rect 21420 16046 21422 16098
rect 21422 16046 21474 16098
rect 21474 16046 21476 16098
rect 21420 16044 21476 16046
rect 21308 15932 21364 15988
rect 19964 15148 20020 15204
rect 20524 15148 20580 15204
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21980 19292 22036 19348
rect 21868 18844 21924 18900
rect 22764 23436 22820 23492
rect 22764 23100 22820 23156
rect 23100 23378 23156 23380
rect 23100 23326 23102 23378
rect 23102 23326 23154 23378
rect 23154 23326 23156 23378
rect 23100 23324 23156 23326
rect 24444 23436 24500 23492
rect 24556 23772 24612 23828
rect 24108 23324 24164 23380
rect 24556 23212 24612 23268
rect 23660 22988 23716 23044
rect 22652 21084 22708 21140
rect 22204 18396 22260 18452
rect 23100 20860 23156 20916
rect 22764 20018 22820 20020
rect 22764 19966 22766 20018
rect 22766 19966 22818 20018
rect 22818 19966 22820 20018
rect 22764 19964 22820 19966
rect 22764 18732 22820 18788
rect 22876 19180 22932 19236
rect 22764 18060 22820 18116
rect 24892 24780 24948 24836
rect 23436 21084 23492 21140
rect 23324 20076 23380 20132
rect 23772 19964 23828 20020
rect 24444 21756 24500 21812
rect 23996 21420 24052 21476
rect 25340 24668 25396 24724
rect 25228 21420 25284 21476
rect 24220 20188 24276 20244
rect 24332 20300 24388 20356
rect 23100 18396 23156 18452
rect 23436 18844 23492 18900
rect 22988 17948 23044 18004
rect 23212 18172 23268 18228
rect 22876 16770 22932 16772
rect 22876 16718 22878 16770
rect 22878 16718 22930 16770
rect 22930 16718 22932 16770
rect 22876 16716 22932 16718
rect 21756 15148 21812 15204
rect 22316 15148 22372 15204
rect 23324 15148 23380 15204
rect 24108 18844 24164 18900
rect 24892 20188 24948 20244
rect 24444 19404 24500 19460
rect 24556 19346 24612 19348
rect 24556 19294 24558 19346
rect 24558 19294 24610 19346
rect 24610 19294 24612 19346
rect 24556 19292 24612 19294
rect 26348 24610 26404 24612
rect 26348 24558 26350 24610
rect 26350 24558 26402 24610
rect 26402 24558 26404 24610
rect 26348 24556 26404 24558
rect 27356 24780 27412 24836
rect 27020 24556 27076 24612
rect 37660 26290 37716 26292
rect 37660 26238 37662 26290
rect 37662 26238 37714 26290
rect 37714 26238 37716 26290
rect 37660 26236 37716 26238
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 39900 25564 39956 25620
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 28364 24668 28420 24724
rect 27020 23826 27076 23828
rect 27020 23774 27022 23826
rect 27022 23774 27074 23826
rect 27074 23774 27076 23826
rect 27020 23772 27076 23774
rect 29484 25282 29540 25284
rect 29484 25230 29486 25282
rect 29486 25230 29538 25282
rect 29538 25230 29540 25282
rect 29484 25228 29540 25230
rect 40012 24892 40068 24948
rect 29260 24668 29316 24724
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 28588 23884 28644 23940
rect 28924 23884 28980 23940
rect 28028 23660 28084 23716
rect 27916 22146 27972 22148
rect 27916 22094 27918 22146
rect 27918 22094 27970 22146
rect 27970 22094 27972 22146
rect 27916 22092 27972 22094
rect 27804 21532 27860 21588
rect 27916 20412 27972 20468
rect 28588 21532 28644 21588
rect 26124 19740 26180 19796
rect 26348 19458 26404 19460
rect 26348 19406 26350 19458
rect 26350 19406 26402 19458
rect 26402 19406 26404 19458
rect 26348 19404 26404 19406
rect 25676 19346 25732 19348
rect 25676 19294 25678 19346
rect 25678 19294 25730 19346
rect 25730 19294 25732 19346
rect 25676 19292 25732 19294
rect 28812 20412 28868 20468
rect 29372 23938 29428 23940
rect 29372 23886 29374 23938
rect 29374 23886 29426 23938
rect 29426 23886 29428 23938
rect 29372 23884 29428 23886
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 29036 23714 29092 23716
rect 29036 23662 29038 23714
rect 29038 23662 29090 23714
rect 29090 23662 29092 23714
rect 29036 23660 29092 23662
rect 29260 23714 29316 23716
rect 29260 23662 29262 23714
rect 29262 23662 29314 23714
rect 29314 23662 29316 23714
rect 29260 23660 29316 23662
rect 30044 23660 30100 23716
rect 40012 23548 40068 23604
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 40012 20860 40068 20916
rect 30044 20412 30100 20468
rect 29708 20130 29764 20132
rect 29708 20078 29710 20130
rect 29710 20078 29762 20130
rect 29762 20078 29764 20130
rect 29708 20076 29764 20078
rect 27244 19516 27300 19572
rect 24892 19180 24948 19236
rect 26684 19234 26740 19236
rect 26684 19182 26686 19234
rect 26686 19182 26738 19234
rect 26738 19182 26740 19234
rect 26684 19180 26740 19182
rect 29372 19516 29428 19572
rect 27804 19234 27860 19236
rect 27804 19182 27806 19234
rect 27806 19182 27858 19234
rect 27858 19182 27860 19234
rect 27804 19180 27860 19182
rect 25228 18732 25284 18788
rect 23548 18450 23604 18452
rect 23548 18398 23550 18450
rect 23550 18398 23602 18450
rect 23602 18398 23604 18450
rect 23548 18396 23604 18398
rect 24332 18562 24388 18564
rect 24332 18510 24334 18562
rect 24334 18510 24386 18562
rect 24386 18510 24388 18562
rect 24332 18508 24388 18510
rect 25116 18508 25172 18564
rect 23884 18396 23940 18452
rect 24332 18226 24388 18228
rect 24332 18174 24334 18226
rect 24334 18174 24386 18226
rect 24386 18174 24388 18226
rect 24332 18172 24388 18174
rect 26460 18956 26516 19012
rect 25900 18338 25956 18340
rect 25900 18286 25902 18338
rect 25902 18286 25954 18338
rect 25954 18286 25956 18338
rect 25900 18284 25956 18286
rect 23660 17948 23716 18004
rect 24556 16828 24612 16884
rect 23884 16770 23940 16772
rect 23884 16718 23886 16770
rect 23886 16718 23938 16770
rect 23938 16718 23940 16770
rect 23884 16716 23940 16718
rect 25340 18226 25396 18228
rect 25340 18174 25342 18226
rect 25342 18174 25394 18226
rect 25394 18174 25396 18226
rect 25340 18172 25396 18174
rect 25340 16882 25396 16884
rect 25340 16830 25342 16882
rect 25342 16830 25394 16882
rect 25394 16830 25396 16882
rect 25340 16828 25396 16830
rect 27356 19010 27412 19012
rect 27356 18958 27358 19010
rect 27358 18958 27410 19010
rect 27410 18958 27412 19010
rect 27356 18956 27412 18958
rect 26572 18338 26628 18340
rect 26572 18286 26574 18338
rect 26574 18286 26626 18338
rect 26626 18286 26628 18338
rect 26572 18284 26628 18286
rect 27468 18396 27524 18452
rect 27692 18508 27748 18564
rect 27020 18284 27076 18340
rect 29260 18508 29316 18564
rect 37660 20076 37716 20132
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 30380 19234 30436 19236
rect 30380 19182 30382 19234
rect 30382 19182 30434 19234
rect 30434 19182 30436 19234
rect 30380 19180 30436 19182
rect 40012 18844 40068 18900
rect 30156 18396 30212 18452
rect 29148 18172 29204 18228
rect 28588 18060 28644 18116
rect 25788 16882 25844 16884
rect 25788 16830 25790 16882
rect 25790 16830 25842 16882
rect 25842 16830 25844 16882
rect 25788 16828 25844 16830
rect 26908 16828 26964 16884
rect 37660 18450 37716 18452
rect 37660 18398 37662 18450
rect 37662 18398 37714 18450
rect 37714 18398 37716 18450
rect 37660 18396 37716 18398
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 30156 18060 30212 18116
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 25228 15538 25284 15540
rect 25228 15486 25230 15538
rect 25230 15486 25282 15538
rect 25282 15486 25284 15538
rect 25228 15484 25284 15486
rect 25900 15538 25956 15540
rect 25900 15486 25902 15538
rect 25902 15486 25954 15538
rect 25954 15486 25956 15538
rect 25900 15484 25956 15486
rect 26348 15484 26404 15540
rect 24556 15202 24612 15204
rect 24556 15150 24558 15202
rect 24558 15150 24610 15202
rect 24610 15150 24612 15202
rect 24556 15148 24612 15150
rect 26236 15426 26292 15428
rect 26236 15374 26238 15426
rect 26238 15374 26290 15426
rect 26290 15374 26292 15426
rect 26236 15372 26292 15374
rect 28588 15372 28644 15428
rect 27020 15260 27076 15316
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19964 4060 20020 4116
rect 20748 4114 20804 4116
rect 20748 4062 20750 4114
rect 20750 4062 20802 4114
rect 20802 4062 20804 4114
rect 20748 4060 20804 4062
rect 21532 3612 21588 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 25564 4060 25620 4116
rect 22428 3666 22484 3668
rect 22428 3614 22430 3666
rect 22430 3614 22482 3666
rect 22482 3614 22484 3666
rect 22428 3612 22484 3614
rect 26796 4114 26852 4116
rect 26796 4062 26798 4114
rect 26798 4062 26850 4114
rect 26850 4062 26852 4114
rect 26796 4060 26852 4062
rect 26236 3612 26292 3668
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 20850 38220 20860 38276
rect 20916 38220 22092 38276
rect 22148 38220 22158 38276
rect 16146 37884 16156 37940
rect 16212 37884 16940 37940
rect 16996 37884 17006 37940
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 17490 37436 17500 37492
rect 17556 37436 18508 37492
rect 18564 37436 18574 37492
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 20850 37212 20860 37268
rect 20916 37212 21644 37268
rect 21700 37212 21710 37268
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 41200 36372 42000 36400
rect 40226 36316 40236 36372
rect 40292 36316 42000 36372
rect 41200 36288 42000 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 0 26292 800 26320
rect 0 26236 4172 26292
rect 4228 26236 4238 26292
rect 27906 26236 27916 26292
rect 27972 26236 37660 26292
rect 37716 26236 37726 26292
rect 0 26208 800 26236
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 41200 25620 42000 25648
rect 16594 25564 16604 25620
rect 16660 25564 17612 25620
rect 17668 25564 18844 25620
rect 18900 25564 18910 25620
rect 39890 25564 39900 25620
rect 39956 25564 42000 25620
rect 41200 25536 42000 25564
rect 4274 25452 4284 25508
rect 4340 25452 11788 25508
rect 11844 25452 11854 25508
rect 31892 25452 37660 25508
rect 37716 25452 37726 25508
rect 31892 25284 31948 25452
rect 13906 25228 13916 25284
rect 13972 25228 14700 25284
rect 14756 25228 17948 25284
rect 18004 25228 19404 25284
rect 19460 25228 19964 25284
rect 20020 25228 20972 25284
rect 21028 25228 21038 25284
rect 29474 25228 29484 25284
rect 29540 25228 31948 25284
rect 13794 25116 13804 25172
rect 13860 25116 15372 25172
rect 15428 25116 15438 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 14802 25004 14812 25060
rect 14868 25004 17724 25060
rect 17780 25004 17790 25060
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 11778 24892 11788 24948
rect 11844 24892 15260 24948
rect 15316 24892 15326 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 18946 24780 18956 24836
rect 19012 24780 20972 24836
rect 21028 24780 24892 24836
rect 24948 24780 27356 24836
rect 27412 24780 27422 24836
rect 15026 24668 15036 24724
rect 15092 24668 17500 24724
rect 17556 24668 17566 24724
rect 17826 24668 17836 24724
rect 17892 24668 18732 24724
rect 18788 24668 19740 24724
rect 19796 24668 19806 24724
rect 21186 24668 21196 24724
rect 21252 24668 23548 24724
rect 23604 24668 24332 24724
rect 24388 24668 25340 24724
rect 25396 24668 25406 24724
rect 28354 24668 28364 24724
rect 28420 24668 29260 24724
rect 29316 24668 37660 24724
rect 37716 24668 37726 24724
rect 26338 24556 26348 24612
rect 26404 24556 27020 24612
rect 27076 24556 27086 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 12674 24220 12684 24276
rect 12740 24220 13468 24276
rect 13524 24220 19516 24276
rect 19572 24220 21196 24276
rect 21252 24220 21262 24276
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 13794 23884 13804 23940
rect 13860 23884 14924 23940
rect 14980 23884 14990 23940
rect 19170 23884 19180 23940
rect 19236 23884 19516 23940
rect 19572 23884 20636 23940
rect 20692 23884 20702 23940
rect 28578 23884 28588 23940
rect 28644 23884 28924 23940
rect 28980 23884 29372 23940
rect 29428 23884 29438 23940
rect 31892 23884 37660 23940
rect 37716 23884 37726 23940
rect 24546 23772 24556 23828
rect 24612 23772 27020 23828
rect 27076 23772 27086 23828
rect 31892 23716 31948 23884
rect 15698 23660 15708 23716
rect 15764 23660 17388 23716
rect 17444 23660 18732 23716
rect 18788 23660 18798 23716
rect 28018 23660 28028 23716
rect 28084 23660 29036 23716
rect 29092 23660 29102 23716
rect 29250 23660 29260 23716
rect 29316 23660 30044 23716
rect 30100 23660 31948 23716
rect 0 23604 800 23632
rect 41200 23604 42000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 14018 23548 14028 23604
rect 14084 23548 17500 23604
rect 17556 23548 19180 23604
rect 19236 23548 19246 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 14924 23492 14980 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 14914 23436 14924 23492
rect 14980 23436 14990 23492
rect 21746 23436 21756 23492
rect 21812 23436 22764 23492
rect 22820 23436 24444 23492
rect 24500 23436 24510 23492
rect 14802 23324 14812 23380
rect 14868 23324 15932 23380
rect 15988 23324 15998 23380
rect 19618 23324 19628 23380
rect 19684 23324 21868 23380
rect 21924 23324 21934 23380
rect 23090 23324 23100 23380
rect 23156 23324 24108 23380
rect 24164 23324 24174 23380
rect 20178 23212 20188 23268
rect 20244 23212 21084 23268
rect 21140 23212 21980 23268
rect 22036 23212 22046 23268
rect 22418 23212 22428 23268
rect 22484 23212 24556 23268
rect 24612 23212 24622 23268
rect 8372 23100 11564 23156
rect 11620 23100 15036 23156
rect 15092 23100 15102 23156
rect 15250 23100 15260 23156
rect 15316 23100 16604 23156
rect 16660 23100 16670 23156
rect 20626 23100 20636 23156
rect 20692 23100 21308 23156
rect 21364 23100 22764 23156
rect 22820 23100 22830 23156
rect 8372 23044 8428 23100
rect 4274 22988 4284 23044
rect 4340 22988 8428 23044
rect 18946 22988 18956 23044
rect 19012 22988 19292 23044
rect 19348 22988 19740 23044
rect 19796 22988 21644 23044
rect 21700 22988 21710 23044
rect 22530 22988 22540 23044
rect 22596 22988 23660 23044
rect 23716 22988 23726 23044
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 1922 22428 1932 22484
rect 1988 22428 1998 22484
rect 0 22260 800 22288
rect 1932 22260 1988 22428
rect 4274 22316 4284 22372
rect 4340 22316 11004 22372
rect 11060 22316 14252 22372
rect 14308 22316 14318 22372
rect 16594 22316 16604 22372
rect 16660 22316 17612 22372
rect 17668 22316 17678 22372
rect 17826 22316 17836 22372
rect 17892 22316 18452 22372
rect 18396 22260 18452 22316
rect 0 22204 1988 22260
rect 12898 22204 12908 22260
rect 12964 22204 14140 22260
rect 14196 22204 14206 22260
rect 15474 22204 15484 22260
rect 15540 22204 16156 22260
rect 16212 22204 16940 22260
rect 16996 22204 18060 22260
rect 18116 22204 18126 22260
rect 18386 22204 18396 22260
rect 18452 22204 18956 22260
rect 19012 22204 19022 22260
rect 19394 22204 19404 22260
rect 19460 22204 22204 22260
rect 22260 22204 22270 22260
rect 0 22176 800 22204
rect 18162 22092 18172 22148
rect 18228 22092 22316 22148
rect 22372 22092 27916 22148
rect 27972 22092 27982 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 17714 21756 17724 21812
rect 17780 21756 18396 21812
rect 18452 21756 18732 21812
rect 18788 21756 18798 21812
rect 21746 21756 21756 21812
rect 21812 21756 24444 21812
rect 24500 21756 24510 21812
rect 17266 21644 17276 21700
rect 17332 21644 19740 21700
rect 19796 21644 19806 21700
rect 20626 21644 20636 21700
rect 20692 21644 22428 21700
rect 22484 21644 22494 21700
rect 17154 21532 17164 21588
rect 17220 21532 18732 21588
rect 18788 21532 19068 21588
rect 19124 21532 19134 21588
rect 19740 21476 19796 21644
rect 20178 21532 20188 21588
rect 20244 21532 21532 21588
rect 21588 21532 21598 21588
rect 27794 21532 27804 21588
rect 27860 21532 28588 21588
rect 28644 21532 37660 21588
rect 37716 21532 37726 21588
rect 19740 21420 23996 21476
rect 24052 21420 25228 21476
rect 25284 21420 25294 21476
rect 18386 21308 18396 21364
rect 18452 21308 19404 21364
rect 19460 21308 20524 21364
rect 20580 21308 20590 21364
rect 18610 21196 18620 21252
rect 18676 21196 19628 21252
rect 19684 21196 19740 21252
rect 19796 21196 19806 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 14578 21084 14588 21140
rect 14644 21084 15932 21140
rect 15988 21084 15998 21140
rect 16706 21084 16716 21140
rect 16772 21084 19964 21140
rect 20020 21084 22428 21140
rect 22484 21084 22494 21140
rect 22642 21084 22652 21140
rect 22708 21084 23436 21140
rect 23492 21084 23502 21140
rect 4162 20972 4172 21028
rect 4228 20972 21308 21028
rect 21364 20972 21374 21028
rect 41200 20916 42000 20944
rect 16482 20860 16492 20916
rect 16548 20860 17556 20916
rect 18274 20860 18284 20916
rect 18340 20860 23100 20916
rect 23156 20860 23166 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 17500 20804 17556 20860
rect 41200 20832 42000 20860
rect 15250 20748 15260 20804
rect 15316 20748 16716 20804
rect 16772 20748 16782 20804
rect 17490 20748 17500 20804
rect 17556 20748 22204 20804
rect 22260 20748 22270 20804
rect 13794 20636 13804 20692
rect 13860 20636 14924 20692
rect 14980 20636 17388 20692
rect 17444 20636 17454 20692
rect 18946 20636 18956 20692
rect 19012 20636 19964 20692
rect 20020 20636 20412 20692
rect 20468 20636 20478 20692
rect 17602 20524 17612 20580
rect 17668 20524 18284 20580
rect 18340 20524 18350 20580
rect 19282 20524 19292 20580
rect 19348 20524 26908 20580
rect 26852 20468 26908 20524
rect 26852 20412 27916 20468
rect 27972 20412 28812 20468
rect 28868 20412 30044 20468
rect 30100 20412 30110 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 22194 20300 22204 20356
rect 22260 20300 24332 20356
rect 24388 20300 24398 20356
rect 0 20244 800 20272
rect 0 20188 1932 20244
rect 1988 20188 1998 20244
rect 14578 20188 14588 20244
rect 14644 20188 16044 20244
rect 16100 20188 17892 20244
rect 18050 20188 18060 20244
rect 18116 20188 22316 20244
rect 22372 20188 24220 20244
rect 24276 20188 24892 20244
rect 24948 20188 24958 20244
rect 0 20160 800 20188
rect 17836 20132 17892 20188
rect 8372 20076 11788 20132
rect 11844 20076 11854 20132
rect 15250 20076 15260 20132
rect 15316 20076 16828 20132
rect 16884 20076 16894 20132
rect 17836 20076 19628 20132
rect 19684 20076 19964 20132
rect 20020 20076 20030 20132
rect 20514 20076 20524 20132
rect 20580 20076 23324 20132
rect 23380 20076 23390 20132
rect 29698 20076 29708 20132
rect 29764 20076 37660 20132
rect 37716 20076 37726 20132
rect 8372 20020 8428 20076
rect 4274 19964 4284 20020
rect 4340 19964 8428 20020
rect 11330 19964 11340 20020
rect 11396 19964 14812 20020
rect 14868 19964 14878 20020
rect 15026 19964 15036 20020
rect 15092 19964 15708 20020
rect 15764 19964 15774 20020
rect 21522 19964 21532 20020
rect 21588 19964 22764 20020
rect 22820 19964 23772 20020
rect 23828 19964 23838 20020
rect 11340 19908 11396 19964
rect 4162 19852 4172 19908
rect 4228 19852 11396 19908
rect 13906 19852 13916 19908
rect 13972 19852 15596 19908
rect 15652 19852 15662 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 19954 19740 19964 19796
rect 20020 19740 26124 19796
rect 26180 19740 26908 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 26852 19572 26908 19740
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 0 19516 1988 19572
rect 26852 19516 27244 19572
rect 27300 19516 29372 19572
rect 29428 19516 29438 19572
rect 0 19488 800 19516
rect 18834 19404 18844 19460
rect 18900 19404 24444 19460
rect 24500 19404 26348 19460
rect 26404 19404 26414 19460
rect 21970 19292 21980 19348
rect 22036 19292 24556 19348
rect 24612 19292 25676 19348
rect 25732 19292 25742 19348
rect 15138 19180 15148 19236
rect 15204 19180 19852 19236
rect 19908 19180 22876 19236
rect 22932 19180 22942 19236
rect 24882 19180 24892 19236
rect 24948 19180 26684 19236
rect 26740 19180 26750 19236
rect 27794 19180 27804 19236
rect 27860 19180 30380 19236
rect 30436 19180 30446 19236
rect 11778 19068 11788 19124
rect 11844 19068 15036 19124
rect 15092 19068 15102 19124
rect 26450 18956 26460 19012
rect 26516 18956 27356 19012
rect 27412 18956 27422 19012
rect 41200 18900 42000 18928
rect 21858 18844 21868 18900
rect 21924 18844 23436 18900
rect 23492 18844 24108 18900
rect 24164 18844 24174 18900
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 22754 18732 22764 18788
rect 22820 18732 25228 18788
rect 25284 18732 25294 18788
rect 24322 18508 24332 18564
rect 24388 18508 25116 18564
rect 25172 18508 25182 18564
rect 27682 18508 27692 18564
rect 27748 18508 29260 18564
rect 29316 18508 29326 18564
rect 16258 18396 16268 18452
rect 16324 18396 17724 18452
rect 17780 18396 18732 18452
rect 18788 18396 19404 18452
rect 19460 18396 19470 18452
rect 22194 18396 22204 18452
rect 22260 18396 23100 18452
rect 23156 18396 23548 18452
rect 23604 18396 23614 18452
rect 23874 18396 23884 18452
rect 23940 18396 27468 18452
rect 27524 18396 27534 18452
rect 30146 18396 30156 18452
rect 30212 18396 37660 18452
rect 37716 18396 37726 18452
rect 23884 18340 23940 18396
rect 19170 18284 19180 18340
rect 19236 18284 19628 18340
rect 19684 18284 23940 18340
rect 25890 18284 25900 18340
rect 25956 18284 26572 18340
rect 26628 18284 27020 18340
rect 27076 18284 27086 18340
rect 41200 18228 42000 18256
rect 23202 18172 23212 18228
rect 23268 18172 24332 18228
rect 24388 18172 24398 18228
rect 25330 18172 25340 18228
rect 25396 18172 29148 18228
rect 29204 18172 29214 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 25340 18116 25396 18172
rect 41200 18144 42000 18172
rect 18946 18060 18956 18116
rect 19012 18060 19740 18116
rect 19796 18060 22764 18116
rect 22820 18060 25396 18116
rect 28578 18060 28588 18116
rect 28644 18060 30156 18116
rect 30212 18060 30222 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 22978 17948 22988 18004
rect 23044 17948 23660 18004
rect 23716 17948 23726 18004
rect 15810 17612 15820 17668
rect 15876 17612 16716 17668
rect 16772 17612 16782 17668
rect 14690 17388 14700 17444
rect 14756 17388 16940 17444
rect 16996 17388 17006 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 4274 16828 4284 16884
rect 4340 16828 13468 16884
rect 13524 16828 13534 16884
rect 14018 16828 14028 16884
rect 14084 16828 16268 16884
rect 16324 16828 16334 16884
rect 16706 16828 16716 16884
rect 16772 16828 18284 16884
rect 18340 16828 18350 16884
rect 24546 16828 24556 16884
rect 24612 16828 25340 16884
rect 25396 16828 25788 16884
rect 25844 16828 26908 16884
rect 26964 16828 26974 16884
rect 17602 16716 17612 16772
rect 17668 16716 18844 16772
rect 18900 16716 18910 16772
rect 22866 16716 22876 16772
rect 22932 16716 23884 16772
rect 23940 16716 23950 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16212 800 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 16258 16156 16268 16212
rect 16324 16156 16604 16212
rect 16660 16156 17052 16212
rect 17108 16156 17500 16212
rect 17556 16156 18956 16212
rect 19012 16156 19022 16212
rect 0 16128 800 16156
rect 18274 16044 18284 16100
rect 18340 16044 19180 16100
rect 19236 16044 19852 16100
rect 19908 16044 19918 16100
rect 20178 16044 20188 16100
rect 20244 16044 21420 16100
rect 21476 16044 21486 16100
rect 19282 15932 19292 15988
rect 19348 15932 20412 15988
rect 20468 15932 21308 15988
rect 21364 15932 21374 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 25218 15484 25228 15540
rect 25284 15484 25900 15540
rect 25956 15484 26348 15540
rect 26404 15484 26414 15540
rect 13458 15372 13468 15428
rect 13524 15372 15596 15428
rect 15652 15372 15662 15428
rect 26012 15316 26068 15484
rect 26226 15372 26236 15428
rect 26292 15372 28588 15428
rect 28644 15372 28654 15428
rect 26012 15260 27020 15316
rect 27076 15260 27086 15316
rect 18946 15148 18956 15204
rect 19012 15148 19964 15204
rect 20020 15148 20524 15204
rect 20580 15148 21756 15204
rect 21812 15148 22316 15204
rect 22372 15148 23324 15204
rect 23380 15148 24556 15204
rect 24612 15148 24622 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 16818 5180 16828 5236
rect 16884 5180 18060 5236
rect 18116 5180 18126 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 19954 4060 19964 4116
rect 20020 4060 20748 4116
rect 20804 4060 20814 4116
rect 25554 4060 25564 4116
rect 25620 4060 26796 4116
rect 26852 4060 26862 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 21522 3612 21532 3668
rect 21588 3612 22428 3668
rect 22484 3612 22494 3668
rect 26226 3612 26236 3668
rect 26292 3612 29372 3668
rect 29428 3612 29438 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 19628 21196 19684 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 19628 20076 19684 20132
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 19628 21252 19684 21262
rect 19628 20132 19684 21196
rect 19628 20066 19684 20076
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _087_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20720 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _088_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _089_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21728 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _090_
timestamp 1698175906
transform 1 0 23408 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _091_
timestamp 1698175906
transform -1 0 23296 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20832 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _093_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _094_
timestamp 1698175906
transform -1 0 22736 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _096_
timestamp 1698175906
transform -1 0 25760 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17472 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _098_
timestamp 1698175906
transform 1 0 21280 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform -1 0 22960 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _100_
timestamp 1698175906
transform 1 0 15008 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15680 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698175906
transform -1 0 23632 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _103_
timestamp 1698175906
transform -1 0 23296 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _106_
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform 1 0 23968 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17472 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _109_
timestamp 1698175906
transform -1 0 19600 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform -1 0 29456 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _111_
timestamp 1698175906
transform -1 0 29568 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _112_
timestamp 1698175906
transform -1 0 28224 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform -1 0 21616 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _114_
timestamp 1698175906
transform -1 0 15344 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 17920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _116_
timestamp 1698175906
transform 1 0 14896 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15344 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_
timestamp 1698175906
transform -1 0 25872 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _120_
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _121_
timestamp 1698175906
transform 1 0 24080 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22624 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _123_
timestamp 1698175906
transform 1 0 23520 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1698175906
transform 1 0 23632 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 25424 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _126_
timestamp 1698175906
transform 1 0 19376 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _127_
timestamp 1698175906
transform 1 0 19936 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23296 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24640 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform 1 0 24304 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform 1 0 19152 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform 1 0 22064 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform -1 0 28224 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform -1 0 27328 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _136_
timestamp 1698175906
transform 1 0 19712 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform 1 0 29456 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _138_
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform -1 0 22064 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _140_
timestamp 1698175906
transform -1 0 20384 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _141_
timestamp 1698175906
transform -1 0 24752 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform -1 0 19152 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19600 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 28672 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 27664 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _146_
timestamp 1698175906
transform -1 0 19488 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _147_
timestamp 1698175906
transform -1 0 19824 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _149_
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20832 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _151_
timestamp 1698175906
transform 1 0 15456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform -1 0 16576 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _153_
timestamp 1698175906
transform -1 0 16464 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _154_
timestamp 1698175906
transform 1 0 16576 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 17808 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _156_
timestamp 1698175906
transform -1 0 17360 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _157_
timestamp 1698175906
transform -1 0 19040 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _158_
timestamp 1698175906
transform -1 0 21056 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _159_
timestamp 1698175906
transform 1 0 21616 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _160_
timestamp 1698175906
transform -1 0 20272 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _161_
timestamp 1698175906
transform 1 0 14448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform -1 0 14224 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform 1 0 29904 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_
timestamp 1698175906
transform 1 0 27104 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _165_
timestamp 1698175906
transform -1 0 15904 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _166_
timestamp 1698175906
transform -1 0 14000 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform 1 0 13888 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform -1 0 13104 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _170_
timestamp 1698175906
transform 1 0 17696 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _171_
timestamp 1698175906
transform -1 0 18256 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform -1 0 28112 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 27104 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14672 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _175_
timestamp 1698175906
transform 1 0 26992 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _176_
timestamp 1698175906
transform -1 0 14896 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23184 0 1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _178_
timestamp 1698175906
transform 1 0 21504 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _179_
timestamp 1698175906
transform 1 0 20384 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _180_
timestamp 1698175906
transform -1 0 25648 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _181_
timestamp 1698175906
transform 1 0 21056 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_
timestamp 1698175906
transform 1 0 25424 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1698175906
transform 1 0 26768 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1698175906
transform -1 0 19712 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1698175906
transform 1 0 26432 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1698175906
transform 1 0 16464 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1698175906
transform 1 0 18816 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1698175906
transform -1 0 16576 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 17696 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform -1 0 14448 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 25536 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform -1 0 14896 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform -1 0 14112 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 13776 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 25536 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _199_
timestamp 1698175906
transform 1 0 25760 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _200_
timestamp 1698175906
transform 1 0 19152 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _201_
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _202_
timestamp 1698175906
transform -1 0 21840 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _203_
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__CLK
timestamp 1698175906
transform 1 0 26768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__CLK
timestamp 1698175906
transform 1 0 26880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__CLK
timestamp 1698175906
transform 1 0 25872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__CLK
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__CLK
timestamp 1698175906
transform 1 0 26320 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__CLK
timestamp 1698175906
transform 1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__CLK
timestamp 1698175906
transform 1 0 25872 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__CLK
timestamp 1698175906
transform 1 0 26544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK
timestamp 1698175906
transform 1 0 19936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__CLK
timestamp 1698175906
transform 1 0 26208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__CLK
timestamp 1698175906
transform 1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__CLK
timestamp 1698175906
transform 1 0 22288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1698175906
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698175906
transform 1 0 14448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 14896 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 14336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 17920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 21168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698175906
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698175906
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_158
timestamp 1698175906
transform 1 0 19040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_162
timestamp 1698175906
transform 1 0 19488 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_189
timestamp 1698175906
transform 1 0 22512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_205
timestamp 1698175906
transform 1 0 24304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 28560 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_173
timestamp 1698175906
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_154
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_185
timestamp 1698175906
transform 1 0 22064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_189
timestamp 1698175906
transform 1 0 22512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_205
timestamp 1698175906
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_131
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_164
timestamp 1698175906
transform 1 0 19712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_168
timestamp 1698175906
transform 1 0 20160 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1698175906
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_130
timestamp 1698175906
transform 1 0 15904 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_158
timestamp 1698175906
transform 1 0 19040 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_165
timestamp 1698175906
transform 1 0 19824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_169
timestamp 1698175906
transform 1 0 20272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_205
timestamp 1698175906
transform 1 0 24304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_224
timestamp 1698175906
transform 1 0 26432 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_256
timestamp 1698175906
transform 1 0 30016 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_272
timestamp 1698175906
transform 1 0 31808 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_142
timestamp 1698175906
transform 1 0 17248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_146
timestamp 1698175906
transform 1 0 17696 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_154
timestamp 1698175906
transform 1 0 18592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_162
timestamp 1698175906
transform 1 0 19488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_183
timestamp 1698175906
transform 1 0 21840 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_191
timestamp 1698175906
transform 1 0 22736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_226
timestamp 1698175906
transform 1 0 26656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_230
timestamp 1698175906
transform 1 0 27104 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_238
timestamp 1698175906
transform 1 0 28000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698175906
transform 1 0 13440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698175906
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_147
timestamp 1698175906
transform 1 0 17808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_149
timestamp 1698175906
transform 1 0 18032 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_160
timestamp 1698175906
transform 1 0 19264 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_164
timestamp 1698175906
transform 1 0 19712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_172
timestamp 1698175906
transform 1 0 20608 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_188
timestamp 1698175906
transform 1 0 22400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_245
timestamp 1698175906
transform 1 0 28784 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_123
timestamp 1698175906
transform 1 0 15120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_143
timestamp 1698175906
transform 1 0 17360 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_159
timestamp 1698175906
transform 1 0 19152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_169
timestamp 1698175906
transform 1 0 20272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_227
timestamp 1698175906
transform 1 0 26768 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_121
timestamp 1698175906
transform 1 0 14896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_125
timestamp 1698175906
transform 1 0 15344 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_133
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698175906
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_148
timestamp 1698175906
transform 1 0 17920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_156
timestamp 1698175906
transform 1 0 18816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_158
timestamp 1698175906
transform 1 0 19040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_165
timestamp 1698175906
transform 1 0 19824 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_217
timestamp 1698175906
transform 1 0 25648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_221
timestamp 1698175906
transform 1 0 26096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_256
timestamp 1698175906
transform 1 0 30016 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_272
timestamp 1698175906
transform 1 0 31808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_125
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_157
timestamp 1698175906
transform 1 0 18928 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_179
timestamp 1698175906
transform 1 0 21392 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_238
timestamp 1698175906
transform 1 0 28000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 28448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_260
timestamp 1698175906
transform 1 0 30464 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_292
timestamp 1698175906
transform 1 0 34048 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 35840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_133
timestamp 1698175906
transform 1 0 16240 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_152
timestamp 1698175906
transform 1 0 18368 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_169
timestamp 1698175906
transform 1 0 20272 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_173
timestamp 1698175906
transform 1 0 20720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_177
timestamp 1698175906
transform 1 0 21168 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_199
timestamp 1698175906
transform 1 0 23632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_201
timestamp 1698175906
transform 1 0 23856 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_256
timestamp 1698175906
transform 1 0 30016 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_272
timestamp 1698175906
transform 1 0 31808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_119
timestamp 1698175906
transform 1 0 14672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_128
timestamp 1698175906
transform 1 0 15680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_144
timestamp 1698175906
transform 1 0 17472 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_154
timestamp 1698175906
transform 1 0 18592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_156
timestamp 1698175906
transform 1 0 18816 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_227
timestamp 1698175906
transform 1 0 26768 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_84
timestamp 1698175906
transform 1 0 10752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_114
timestamp 1698175906
transform 1 0 14112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_118
timestamp 1698175906
transform 1 0 14560 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_174
timestamp 1698175906
transform 1 0 20832 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_178
timestamp 1698175906
transform 1 0 21280 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_218
timestamp 1698175906
transform 1 0 25760 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_239
timestamp 1698175906
transform 1 0 28112 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_271
timestamp 1698175906
transform 1 0 31696 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_85
timestamp 1698175906
transform 1 0 10864 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_93
timestamp 1698175906
transform 1 0 11760 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_97
timestamp 1698175906
transform 1 0 12208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_120
timestamp 1698175906
transform 1 0 14784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_128
timestamp 1698175906
transform 1 0 15680 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_136
timestamp 1698175906
transform 1 0 16576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_158
timestamp 1698175906
transform 1 0 19040 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_190
timestamp 1698175906
transform 1 0 22624 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_194
timestamp 1698175906
transform 1 0 23072 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_208
timestamp 1698175906
transform 1 0 24640 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_224
timestamp 1698175906
transform 1 0 26432 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_232
timestamp 1698175906
transform 1 0 27328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_234
timestamp 1698175906
transform 1 0 27552 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_240
timestamp 1698175906
transform 1 0 28224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_128
timestamp 1698175906
transform 1 0 15680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_132
timestamp 1698175906
transform 1 0 16128 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_158
timestamp 1698175906
transform 1 0 19040 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_162
timestamp 1698175906
transform 1 0 19488 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_189
timestamp 1698175906
transform 1 0 22512 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698175906
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_224
timestamp 1698175906
transform 1 0 26432 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_226
timestamp 1698175906
transform 1 0 26656 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_258
timestamp 1698175906
transform 1 0 30240 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698175906
transform 1 0 32032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_113
timestamp 1698175906
transform 1 0 14000 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_123
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_139
timestamp 1698175906
transform 1 0 16912 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_147
timestamp 1698175906
transform 1 0 17808 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_151
timestamp 1698175906
transform 1 0 18256 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_232
timestamp 1698175906
transform 1 0 27328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_236
timestamp 1698175906
transform 1 0 27776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_238
timestamp 1698175906
transform 1 0 28000 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_252
timestamp 1698175906
transform 1 0 29568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_284
timestamp 1698175906
transform 1 0 33152 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_300
timestamp 1698175906
transform 1 0 34944 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_308
timestamp 1698175906
transform 1 0 35840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698175906
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698175906
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698175906
transform 1 0 15904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_151
timestamp 1698175906
transform 1 0 18256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_153
timestamp 1698175906
transform 1 0 18480 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_214
timestamp 1698175906
transform 1 0 25312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_244
timestamp 1698175906
transform 1 0 28672 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_113
timestamp 1698175906
transform 1 0 14000 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_129
timestamp 1698175906
transform 1 0 15792 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_133
timestamp 1698175906
transform 1 0 16240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_164
timestamp 1698175906
transform 1 0 19712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698175906
transform 1 0 20160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698175906
transform 1 0 22064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_187
timestamp 1698175906
transform 1 0 22288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_217
timestamp 1698175906
transform 1 0 25648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_221
timestamp 1698175906
transform 1 0 26096 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_225
timestamp 1698175906
transform 1 0 26544 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_229
timestamp 1698175906
transform 1 0 26992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698175906
transform 1 0 28224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_253
timestamp 1698175906
transform 1 0 29680 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_285
timestamp 1698175906
transform 1 0 33264 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_301
timestamp 1698175906
transform 1 0 35056 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698175906
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698175906
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 13440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 13664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_150
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_166
timestamp 1698175906
transform 1 0 19936 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_174
timestamp 1698175906
transform 1 0 20832 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_177
timestamp 1698175906
transform 1 0 21168 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_193
timestamp 1698175906
transform 1 0 22960 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_201
timestamp 1698175906
transform 1 0 23856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698175906
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_253
timestamp 1698175906
transform 1 0 29680 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_269
timestamp 1698175906
transform 1 0 31472 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_139
timestamp 1698175906
transform 1 0 16912 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_143
timestamp 1698175906
transform 1 0 17360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_145
timestamp 1698175906
transform 1 0 17584 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_183
timestamp 1698175906
transform 1 0 21840 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_215
timestamp 1698175906
transform 1 0 25424 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_231
timestamp 1698175906
transform 1 0 27216 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698175906
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698175906
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_341
timestamp 1698175906
transform 1 0 39536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 23856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 24080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_206
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita64_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17248 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita64_26
timestamp 1698175906
transform 1 0 39984 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 17360 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 16912 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 27328 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 19600 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 25648 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 36288 42000 36400 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 26488 17976 26488 17976 0 _000_
rlabel metal2 13944 24864 13944 24864 0 _001_
rlabel metal2 13160 21728 13160 21728 0 _002_
rlabel metal2 14840 25592 14840 25592 0 _003_
rlabel metal2 26600 19600 26600 19600 0 _004_
rlabel metal2 13664 23240 13664 23240 0 _005_
rlabel metal2 27944 22792 27944 22792 0 _006_
rlabel metal2 13944 19152 13944 19152 0 _007_
rlabel metal2 24136 15736 24136 15736 0 _008_
rlabel metal2 22400 19320 22400 19320 0 _009_
rlabel metal2 20664 16128 20664 16128 0 _010_
rlabel metal2 24752 24920 24752 24920 0 _011_
rlabel metal2 22288 22568 22288 22568 0 _012_
rlabel metal2 27048 24360 27048 24360 0 _013_
rlabel metal2 27720 18480 27720 18480 0 _014_
rlabel metal2 18704 25368 18704 25368 0 _015_
rlabel metal2 27384 25928 27384 25928 0 _016_
rlabel metal3 18256 16744 18256 16744 0 _017_
rlabel metal2 19992 15512 19992 15512 0 _018_
rlabel metal2 15624 16800 15624 16800 0 _019_
rlabel metal2 14728 17192 14728 17192 0 _020_
rlabel metal2 18648 26908 18648 26908 0 _021_
rlabel metal2 13720 19656 13720 19656 0 _022_
rlabel metal3 19936 23912 19936 23912 0 _023_
rlabel metal2 27384 25032 27384 25032 0 _024_
rlabel metal2 19432 24192 19432 24192 0 _025_
rlabel metal2 28168 24192 28168 24192 0 _026_
rlabel metal2 19096 16296 19096 16296 0 _027_
rlabel metal2 18312 16352 18312 16352 0 _028_
rlabel metal3 20832 16072 20832 16072 0 _029_
rlabel metal2 15848 15512 15848 15512 0 _030_
rlabel metal2 14616 21672 14616 21672 0 _031_
rlabel metal2 16856 19096 16856 19096 0 _032_
rlabel metal2 17304 17304 17304 17304 0 _033_
rlabel metal3 18816 24696 18816 24696 0 _034_
rlabel metal2 20216 24696 20216 24696 0 _035_
rlabel metal3 20776 23352 20776 23352 0 _036_
rlabel metal2 14168 19432 14168 19432 0 _037_
rlabel metal3 29120 19208 29120 19208 0 _038_
rlabel metal2 13832 25256 13832 25256 0 _039_
rlabel metal3 13552 22232 13552 22232 0 _040_
rlabel metal2 17584 24920 17584 24920 0 _041_
rlabel metal2 17920 20888 17920 20888 0 _042_
rlabel metal2 27608 20860 27608 20860 0 _043_
rlabel metal2 19992 20720 19992 20720 0 _044_
rlabel metal2 17192 21112 17192 21112 0 _045_
rlabel metal2 22232 19208 22232 19208 0 _046_
rlabel metal2 27496 18704 27496 18704 0 _047_
rlabel metal3 21000 23128 21000 23128 0 _048_
rlabel metal2 19432 21168 19432 21168 0 _049_
rlabel metal2 14952 23408 14952 23408 0 _050_
rlabel metal2 22232 21000 22232 21000 0 _051_
rlabel metal2 16632 22456 16632 22456 0 _052_
rlabel metal2 17304 21336 17304 21336 0 _053_
rlabel metal3 17528 22232 17528 22232 0 _054_
rlabel metal2 22792 19376 22792 19376 0 _055_
rlabel metal2 19992 21336 19992 21336 0 _056_
rlabel metal2 15512 23968 15512 23968 0 _057_
rlabel metal2 15064 23632 15064 23632 0 _058_
rlabel metal3 17976 20552 17976 20552 0 _059_
rlabel metal2 21784 23408 21784 23408 0 _060_
rlabel metal3 19544 23016 19544 23016 0 _061_
rlabel metal2 13496 24192 13496 24192 0 _062_
rlabel metal2 24472 19768 24472 19768 0 _063_
rlabel metal3 20272 22120 20272 22120 0 _064_
rlabel metal3 29456 20440 29456 20440 0 _065_
rlabel metal2 28560 23912 28560 23912 0 _066_
rlabel metal2 28056 23016 28056 23016 0 _067_
rlabel metal2 19880 19600 19880 19600 0 _068_
rlabel metal2 15064 19712 15064 19712 0 _069_
rlabel metal2 14952 20720 14952 20720 0 _070_
rlabel metal2 15568 20104 15568 20104 0 _071_
rlabel metal2 16072 20160 16072 20160 0 _072_
rlabel metal2 25424 18984 25424 18984 0 _073_
rlabel metal2 29176 18592 29176 18592 0 _074_
rlabel metal2 23240 17640 23240 17640 0 _075_
rlabel metal3 23408 16744 23408 16744 0 _076_
rlabel metal2 23968 15288 23968 15288 0 _077_
rlabel metal2 20216 17136 20216 17136 0 _078_
rlabel metal2 24304 22344 24304 22344 0 _079_
rlabel metal2 24584 24304 24584 24304 0 _080_
rlabel metal2 17752 18480 17752 18480 0 _081_
rlabel metal2 19656 20832 19656 20832 0 _082_
rlabel metal2 27160 24136 27160 24136 0 _083_
rlabel metal2 27272 19376 27272 19376 0 _084_
rlabel metal2 29736 19488 29736 19488 0 _085_
rlabel metal3 20888 21560 20888 21560 0 _086_
rlabel metal3 2478 26264 2478 26264 0 clk
rlabel metal2 23576 21000 23576 21000 0 clknet_0_clk
rlabel metal2 26936 16520 26936 16520 0 clknet_1_0__leaf_clk
rlabel metal2 27160 23240 27160 23240 0 clknet_1_1__leaf_clk
rlabel metal2 25760 19320 25760 19320 0 dut64.count\[0\]
rlabel metal2 24248 19432 24248 19432 0 dut64.count\[1\]
rlabel metal2 23688 22792 23688 22792 0 dut64.count\[2\]
rlabel metal2 24136 23856 24136 23856 0 dut64.count\[3\]
rlabel metal2 28616 9464 28616 9464 0 net1
rlabel metal2 13496 16520 13496 16520 0 net10
rlabel metal2 19600 14392 19600 14392 0 net11
rlabel metal2 19320 15568 19320 15568 0 net12
rlabel metal3 30716 25256 30716 25256 0 net13
rlabel metal2 4200 20328 4200 20328 0 net14
rlabel metal2 30184 18536 30184 18536 0 net15
rlabel metal3 17752 25592 17752 25592 0 net16
rlabel metal2 21336 32480 21336 32480 0 net17
rlabel metal2 27944 25816 27944 25816 0 net18
rlabel metal2 25592 15260 25592 15260 0 net19
rlabel metal2 29288 25088 29288 25088 0 net2
rlabel metal3 6356 19992 6356 19992 0 net20
rlabel metal2 4312 23464 4312 23464 0 net21
rlabel metal2 30072 23352 30072 23352 0 net22
rlabel metal2 29848 19208 29848 19208 0 net23
rlabel metal2 27832 21616 27832 21616 0 net24
rlabel metal3 16576 37912 16576 37912 0 net25
rlabel metal3 40754 36344 40754 36344 0 net26
rlabel metal2 11032 21896 11032 21896 0 net3
rlabel metal2 17472 31920 17472 31920 0 net4
rlabel metal2 17528 16856 17528 16856 0 net5
rlabel metal2 27048 9408 27048 9408 0 net6
rlabel metal2 11816 25032 11816 25032 0 net7
rlabel metal3 21280 37240 21280 37240 0 net8
rlabel metal2 21840 13608 21840 13608 0 net9
rlabel metal2 26264 2198 26264 2198 0 segm[0]
rlabel metal2 40040 24360 40040 24360 0 segm[10]
rlabel metal3 1358 22232 1358 22232 0 segm[11]
rlabel metal2 17528 39354 17528 39354 0 segm[12]
rlabel metal3 17472 5208 17472 5208 0 segm[13]
rlabel metal2 24248 2058 24248 2058 0 segm[2]
rlabel metal3 1358 24920 1358 24920 0 segm[3]
rlabel metal2 20216 39354 20216 39354 0 segm[5]
rlabel metal3 22008 3640 22008 3640 0 segm[6]
rlabel metal3 1358 16184 1358 16184 0 segm[7]
rlabel metal2 19544 2058 19544 2058 0 segm[8]
rlabel metal2 18872 2198 18872 2198 0 segm[9]
rlabel metal2 40040 25256 40040 25256 0 sel[0]
rlabel metal3 1358 20216 1358 20216 0 sel[10]
rlabel metal3 40642 18200 40642 18200 0 sel[11]
rlabel metal2 19544 39746 19544 39746 0 sel[1]
rlabel metal2 20888 39746 20888 39746 0 sel[2]
rlabel metal2 39928 25872 39928 25872 0 sel[3]
rlabel metal3 26208 4088 26208 4088 0 sel[4]
rlabel metal3 1358 19544 1358 19544 0 sel[5]
rlabel metal3 1358 23576 1358 23576 0 sel[6]
rlabel metal2 40040 23800 40040 23800 0 sel[7]
rlabel metal2 40040 19096 40040 19096 0 sel[8]
rlabel metal2 40040 21112 40040 21112 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
