magic
tech gf180mcuD
magscale 1 5
timestamp 1699641544
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9031 19137 9057 19143
rect 9031 19105 9057 19111
rect 11047 19137 11073 19143
rect 11047 19105 11073 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 14687 19137 14713 19143
rect 14687 19105 14713 19111
rect 8521 18999 8527 19025
rect 8553 18999 8559 19025
rect 10537 18999 10543 19025
rect 10569 18999 10575 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 14289 18999 14295 19025
rect 14321 18999 14327 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10711 18745 10737 18751
rect 10711 18713 10737 18719
rect 13399 18745 13425 18751
rect 13399 18713 13425 18719
rect 10201 18607 10207 18633
rect 10233 18607 10239 18633
rect 13113 18607 13119 18633
rect 13145 18607 13151 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 967 13593 993 13599
rect 20007 13593 20033 13599
rect 8521 13567 8527 13593
rect 8553 13567 8559 13593
rect 10369 13567 10375 13593
rect 10401 13567 10407 13593
rect 13169 13567 13175 13593
rect 13201 13567 13207 13593
rect 967 13561 993 13567
rect 20007 13561 20033 13567
rect 2137 13511 2143 13537
rect 2169 13511 2175 13537
rect 7065 13511 7071 13537
rect 7097 13511 7103 13537
rect 8913 13511 8919 13537
rect 8945 13511 8951 13537
rect 11769 13511 11775 13537
rect 11801 13511 11807 13537
rect 18937 13511 18943 13537
rect 18969 13511 18975 13537
rect 13399 13481 13425 13487
rect 7457 13455 7463 13481
rect 7489 13455 7495 13481
rect 9305 13455 9311 13481
rect 9337 13455 9343 13481
rect 12105 13455 12111 13481
rect 12137 13455 12143 13481
rect 13399 13449 13425 13455
rect 8751 13425 8777 13431
rect 8751 13393 8777 13399
rect 10711 13425 10737 13431
rect 10711 13393 10737 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7855 13257 7881 13263
rect 7855 13225 7881 13231
rect 12671 13257 12697 13263
rect 13113 13231 13119 13257
rect 13145 13231 13151 13257
rect 12671 13225 12697 13231
rect 8247 13201 8273 13207
rect 8247 13169 8273 13175
rect 10431 13201 10457 13207
rect 10431 13169 10457 13175
rect 12727 13201 12753 13207
rect 12727 13169 12753 13175
rect 8023 13145 8049 13151
rect 7457 13119 7463 13145
rect 7489 13119 7495 13145
rect 7737 13119 7743 13145
rect 7769 13119 7775 13145
rect 8023 13113 8049 13119
rect 8359 13145 8385 13151
rect 12335 13145 12361 13151
rect 8745 13119 8751 13145
rect 8777 13119 8783 13145
rect 10705 13119 10711 13145
rect 10737 13119 10743 13145
rect 8359 13113 8385 13119
rect 12335 13113 12361 13119
rect 12951 13145 12977 13151
rect 13449 13119 13455 13145
rect 13481 13119 13487 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 12951 13113 12977 13119
rect 8135 13089 8161 13095
rect 15079 13089 15105 13095
rect 6057 13063 6063 13089
rect 6089 13063 6095 13089
rect 7121 13063 7127 13089
rect 7153 13063 7159 13089
rect 9137 13063 9143 13089
rect 9169 13063 9175 13089
rect 10201 13063 10207 13089
rect 10233 13063 10239 13089
rect 11041 13063 11047 13089
rect 11073 13063 11079 13089
rect 12105 13063 12111 13089
rect 12137 13063 12143 13089
rect 13785 13063 13791 13089
rect 13817 13063 13823 13089
rect 14849 13063 14855 13089
rect 14881 13063 14887 13089
rect 8135 13057 8161 13063
rect 15079 13057 15105 13063
rect 7911 13033 7937 13039
rect 7911 13001 7937 13007
rect 12615 13033 12641 13039
rect 12615 13001 12641 13007
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 7015 12865 7041 12871
rect 7015 12833 7041 12839
rect 10263 12865 10289 12871
rect 10263 12833 10289 12839
rect 11551 12865 11577 12871
rect 13735 12865 13761 12871
rect 12609 12839 12615 12865
rect 12641 12839 12647 12865
rect 11551 12833 11577 12839
rect 13735 12833 13761 12839
rect 967 12809 993 12815
rect 967 12777 993 12783
rect 10711 12809 10737 12815
rect 10711 12777 10737 12783
rect 11271 12809 11297 12815
rect 11271 12777 11297 12783
rect 10039 12753 10065 12759
rect 11103 12753 11129 12759
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 7849 12727 7855 12753
rect 7881 12727 7887 12753
rect 9697 12727 9703 12753
rect 9729 12727 9735 12753
rect 10089 12727 10095 12753
rect 10121 12727 10127 12753
rect 10039 12721 10065 12727
rect 11103 12721 11129 12727
rect 11383 12753 11409 12759
rect 11383 12721 11409 12727
rect 12335 12753 12361 12759
rect 12335 12721 12361 12727
rect 14295 12753 14321 12759
rect 14295 12721 14321 12727
rect 14799 12753 14825 12759
rect 14799 12721 14825 12727
rect 6959 12697 6985 12703
rect 6959 12665 6985 12671
rect 7519 12697 7545 12703
rect 7519 12665 7545 12671
rect 7575 12697 7601 12703
rect 7575 12665 7601 12671
rect 7631 12697 7657 12703
rect 7631 12665 7657 12671
rect 9535 12697 9561 12703
rect 9535 12665 9561 12671
rect 9983 12697 10009 12703
rect 9983 12665 10009 12671
rect 10655 12697 10681 12703
rect 10655 12665 10681 12671
rect 11159 12697 11185 12703
rect 11159 12665 11185 12671
rect 11495 12697 11521 12703
rect 11495 12665 11521 12671
rect 11551 12697 11577 12703
rect 11551 12665 11577 12671
rect 12279 12697 12305 12703
rect 12279 12665 12305 12671
rect 12391 12697 12417 12703
rect 12391 12665 12417 12671
rect 12783 12697 12809 12703
rect 12783 12665 12809 12671
rect 12839 12697 12865 12703
rect 12839 12665 12865 12671
rect 12951 12697 12977 12703
rect 12951 12665 12977 12671
rect 13791 12697 13817 12703
rect 13791 12665 13817 12671
rect 14239 12697 14265 12703
rect 14239 12665 14265 12671
rect 14519 12697 14545 12703
rect 14519 12665 14545 12671
rect 14631 12697 14657 12703
rect 14631 12665 14657 12671
rect 14687 12697 14713 12703
rect 14687 12665 14713 12671
rect 14911 12697 14937 12703
rect 14911 12665 14937 12671
rect 14967 12697 14993 12703
rect 14967 12665 14993 12671
rect 7239 12641 7265 12647
rect 7239 12609 7265 12615
rect 7463 12641 7489 12647
rect 7463 12609 7489 12615
rect 8079 12641 8105 12647
rect 8079 12609 8105 12615
rect 9591 12641 9617 12647
rect 9591 12609 9617 12615
rect 9927 12641 9953 12647
rect 9927 12609 9953 12615
rect 10767 12641 10793 12647
rect 10767 12609 10793 12615
rect 13735 12641 13761 12647
rect 13735 12609 13761 12615
rect 14127 12641 14153 12647
rect 14127 12609 14153 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7351 12473 7377 12479
rect 7351 12441 7377 12447
rect 9759 12473 9785 12479
rect 9759 12441 9785 12447
rect 13679 12473 13705 12479
rect 13679 12441 13705 12447
rect 10263 12417 10289 12423
rect 6673 12391 6679 12417
rect 6705 12391 6711 12417
rect 14233 12391 14239 12417
rect 14265 12391 14271 12417
rect 10263 12385 10289 12391
rect 7295 12361 7321 12367
rect 8639 12361 8665 12367
rect 7065 12335 7071 12361
rect 7097 12335 7103 12361
rect 7401 12335 7407 12361
rect 7433 12335 7439 12361
rect 7681 12335 7687 12361
rect 7713 12335 7719 12361
rect 7295 12329 7321 12335
rect 8639 12329 8665 12335
rect 8863 12361 8889 12367
rect 8863 12329 8889 12335
rect 8975 12361 9001 12367
rect 10207 12361 10233 12367
rect 9641 12335 9647 12361
rect 9673 12335 9679 12361
rect 9977 12335 9983 12361
rect 10009 12335 10015 12361
rect 13841 12335 13847 12361
rect 13873 12335 13879 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 8975 12329 9001 12335
rect 10207 12329 10233 12335
rect 8919 12305 8945 12311
rect 5609 12279 5615 12305
rect 5641 12279 5647 12305
rect 15297 12279 15303 12305
rect 15329 12279 15335 12305
rect 8919 12273 8945 12279
rect 9815 12249 9841 12255
rect 7569 12223 7575 12249
rect 7601 12223 7607 12249
rect 9815 12217 9841 12223
rect 10095 12249 10121 12255
rect 10095 12217 10121 12223
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 7183 12081 7209 12087
rect 7183 12049 7209 12055
rect 11103 12081 11129 12087
rect 11103 12049 11129 12055
rect 7127 12025 7153 12031
rect 10767 12025 10793 12031
rect 9529 11999 9535 12025
rect 9561 11999 9567 12025
rect 7127 11993 7153 11999
rect 10767 11993 10793 11999
rect 14295 12025 14321 12031
rect 16025 11999 16031 12025
rect 16057 11999 16063 12025
rect 14295 11993 14321 11999
rect 9255 11969 9281 11975
rect 11047 11969 11073 11975
rect 9361 11943 9367 11969
rect 9393 11943 9399 11969
rect 9255 11937 9281 11943
rect 11047 11937 11073 11943
rect 11439 11969 11465 11975
rect 14569 11943 14575 11969
rect 14601 11943 14607 11969
rect 11439 11937 11465 11943
rect 9815 11913 9841 11919
rect 8353 11887 8359 11913
rect 8385 11887 8391 11913
rect 9815 11881 9841 11887
rect 9871 11913 9897 11919
rect 14961 11887 14967 11913
rect 14993 11887 14999 11913
rect 9871 11881 9897 11887
rect 7407 11857 7433 11863
rect 7407 11825 7433 11831
rect 8527 11857 8553 11863
rect 9983 11857 10009 11863
rect 9025 11831 9031 11857
rect 9057 11831 9063 11857
rect 8527 11825 8553 11831
rect 9983 11825 10009 11831
rect 10711 11857 10737 11863
rect 10711 11825 10737 11831
rect 10823 11857 10849 11863
rect 10823 11825 10849 11831
rect 11159 11857 11185 11863
rect 11159 11825 11185 11831
rect 11271 11857 11297 11863
rect 11271 11825 11297 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 8863 11689 8889 11695
rect 7793 11663 7799 11689
rect 7825 11663 7831 11689
rect 8863 11657 8889 11663
rect 9367 11689 9393 11695
rect 9367 11657 9393 11663
rect 10431 11689 10457 11695
rect 10431 11657 10457 11663
rect 10655 11689 10681 11695
rect 11775 11689 11801 11695
rect 11153 11663 11159 11689
rect 11185 11663 11191 11689
rect 10655 11657 10681 11663
rect 11775 11657 11801 11663
rect 12783 11689 12809 11695
rect 12783 11657 12809 11663
rect 14687 11689 14713 11695
rect 14687 11657 14713 11663
rect 14799 11689 14825 11695
rect 14799 11657 14825 11663
rect 15191 11689 15217 11695
rect 15191 11657 15217 11663
rect 8807 11633 8833 11639
rect 8807 11601 8833 11607
rect 8975 11633 9001 11639
rect 8975 11601 9001 11607
rect 9087 11633 9113 11639
rect 9815 11633 9841 11639
rect 9529 11607 9535 11633
rect 9561 11607 9567 11633
rect 9087 11601 9113 11607
rect 9815 11601 9841 11607
rect 10319 11633 10345 11639
rect 10319 11601 10345 11607
rect 10543 11633 10569 11639
rect 10543 11601 10569 11607
rect 11831 11633 11857 11639
rect 11831 11601 11857 11607
rect 13343 11633 13369 11639
rect 13343 11601 13369 11607
rect 7351 11577 7377 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 7065 11551 7071 11577
rect 7097 11551 7103 11577
rect 7351 11545 7377 11551
rect 7519 11577 7545 11583
rect 7519 11545 7545 11551
rect 7631 11577 7657 11583
rect 7631 11545 7657 11551
rect 7967 11577 7993 11583
rect 7967 11545 7993 11551
rect 10263 11577 10289 11583
rect 10991 11577 11017 11583
rect 10761 11551 10767 11577
rect 10793 11551 10799 11577
rect 10263 11545 10289 11551
rect 10991 11545 11017 11551
rect 11663 11577 11689 11583
rect 11663 11545 11689 11551
rect 12671 11577 12697 11583
rect 12671 11545 12697 11551
rect 13007 11577 13033 11583
rect 13007 11545 13033 11551
rect 13231 11577 13257 11583
rect 13231 11545 13257 11551
rect 13399 11577 13425 11583
rect 13399 11545 13425 11551
rect 14855 11577 14881 11583
rect 14855 11545 14881 11551
rect 15079 11577 15105 11583
rect 15079 11545 15105 11551
rect 15247 11577 15273 11583
rect 15247 11545 15273 11551
rect 7407 11521 7433 11527
rect 5609 11495 5615 11521
rect 5641 11495 5647 11521
rect 6673 11495 6679 11521
rect 6705 11495 6711 11521
rect 7407 11489 7433 11495
rect 9759 11521 9785 11527
rect 12727 11521 12753 11527
rect 10649 11495 10655 11521
rect 10681 11495 10687 11521
rect 9759 11489 9785 11495
rect 12727 11489 12753 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 9703 11465 9729 11471
rect 9703 11433 9729 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 7183 11297 7209 11303
rect 7183 11265 7209 11271
rect 14015 11241 14041 11247
rect 9193 11215 9199 11241
rect 9225 11215 9231 11241
rect 12721 11215 12727 11241
rect 12753 11215 12759 11241
rect 13785 11215 13791 11241
rect 13817 11215 13823 11241
rect 14015 11209 14041 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7239 11185 7265 11191
rect 7239 11153 7265 11159
rect 7855 11185 7881 11191
rect 10767 11185 10793 11191
rect 7905 11159 7911 11185
rect 7937 11159 7943 11185
rect 9529 11159 9535 11185
rect 9561 11159 9567 11185
rect 9697 11159 9703 11185
rect 9729 11159 9735 11185
rect 7855 11153 7881 11159
rect 10767 11153 10793 11159
rect 11047 11185 11073 11191
rect 11047 11153 11073 11159
rect 11103 11185 11129 11191
rect 11103 11153 11129 11159
rect 11327 11185 11353 11191
rect 11327 11153 11353 11159
rect 11999 11185 12025 11191
rect 12385 11159 12391 11185
rect 12417 11159 12423 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 11999 11153 12025 11159
rect 7183 11129 7209 11135
rect 7183 11097 7209 11103
rect 7631 11129 7657 11135
rect 10991 11129 11017 11135
rect 7737 11103 7743 11129
rect 7769 11103 7775 11129
rect 9473 11103 9479 11129
rect 9505 11103 9511 11129
rect 9977 11103 9983 11129
rect 10009 11103 10015 11129
rect 7631 11097 7657 11103
rect 10991 11097 11017 11103
rect 11495 11129 11521 11135
rect 11495 11097 11521 11103
rect 12055 11129 12081 11135
rect 12055 11097 12081 11103
rect 7687 11073 7713 11079
rect 7687 11041 7713 11047
rect 10655 11073 10681 11079
rect 10655 11041 10681 11047
rect 12167 11073 12193 11079
rect 12167 11041 12193 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 14911 10905 14937 10911
rect 8409 10879 8415 10905
rect 8441 10879 8447 10905
rect 11937 10879 11943 10905
rect 11969 10879 11975 10905
rect 14911 10873 14937 10879
rect 11551 10849 11577 10855
rect 6057 10823 6063 10849
rect 6089 10823 6095 10849
rect 9249 10823 9255 10849
rect 9281 10823 9287 10849
rect 14681 10823 14687 10849
rect 14713 10823 14719 10849
rect 11551 10817 11577 10823
rect 11495 10793 11521 10799
rect 5665 10767 5671 10793
rect 5697 10767 5703 10793
rect 8297 10767 8303 10793
rect 8329 10767 8335 10793
rect 11321 10767 11327 10793
rect 11353 10767 11359 10793
rect 11495 10761 11521 10767
rect 11663 10793 11689 10799
rect 11663 10761 11689 10767
rect 12111 10793 12137 10799
rect 14519 10793 14545 10799
rect 12889 10767 12895 10793
rect 12921 10767 12927 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 12111 10761 12137 10767
rect 14519 10761 14545 10767
rect 7351 10737 7377 10743
rect 20007 10737 20033 10743
rect 7121 10711 7127 10737
rect 7153 10711 7159 10737
rect 13281 10711 13287 10737
rect 13313 10711 13319 10737
rect 14345 10711 14351 10737
rect 14377 10711 14383 10737
rect 7351 10705 7377 10711
rect 20007 10705 20033 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7519 10513 7545 10519
rect 7519 10481 7545 10487
rect 10039 10513 10065 10519
rect 10039 10481 10065 10487
rect 10319 10513 10345 10519
rect 10319 10481 10345 10487
rect 10655 10513 10681 10519
rect 10655 10481 10681 10487
rect 7967 10457 7993 10463
rect 7967 10425 7993 10431
rect 9479 10457 9505 10463
rect 9479 10425 9505 10431
rect 10935 10457 10961 10463
rect 20007 10457 20033 10463
rect 12889 10431 12895 10457
rect 12921 10431 12927 10457
rect 16081 10431 16087 10457
rect 16113 10431 16119 10457
rect 10935 10425 10961 10431
rect 20007 10425 20033 10431
rect 7463 10401 7489 10407
rect 8527 10401 8553 10407
rect 8241 10375 8247 10401
rect 8273 10375 8279 10401
rect 7463 10369 7489 10375
rect 8527 10369 8553 10375
rect 8639 10401 8665 10407
rect 8639 10369 8665 10375
rect 8807 10401 8833 10407
rect 10823 10401 10849 10407
rect 9249 10375 9255 10401
rect 9281 10375 9287 10401
rect 9753 10375 9759 10401
rect 9785 10375 9791 10401
rect 10369 10375 10375 10401
rect 10401 10375 10407 10401
rect 8807 10369 8833 10375
rect 10823 10369 10849 10375
rect 11103 10401 11129 10407
rect 11209 10375 11215 10401
rect 11241 10375 11247 10401
rect 11657 10375 11663 10401
rect 11689 10375 11695 10401
rect 14625 10375 14631 10401
rect 14657 10375 14663 10401
rect 16305 10375 16311 10401
rect 16337 10375 16343 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 11103 10369 11129 10375
rect 9983 10345 10009 10351
rect 8353 10319 8359 10345
rect 8385 10319 8391 10345
rect 9983 10313 10009 10319
rect 10151 10345 10177 10351
rect 16423 10345 16449 10351
rect 15017 10319 15023 10345
rect 15049 10319 15055 10345
rect 10151 10313 10177 10319
rect 16423 10313 16449 10319
rect 7687 10289 7713 10295
rect 7687 10257 7713 10263
rect 8583 10289 8609 10295
rect 8583 10257 8609 10263
rect 9871 10289 9897 10295
rect 9871 10257 9897 10263
rect 10263 10289 10289 10295
rect 10263 10257 10289 10263
rect 11159 10289 11185 10295
rect 11159 10257 11185 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 8079 10121 8105 10127
rect 9031 10121 9057 10127
rect 8241 10095 8247 10121
rect 8273 10095 8279 10121
rect 8079 10089 8105 10095
rect 9031 10089 9057 10095
rect 13119 10121 13145 10127
rect 13119 10089 13145 10095
rect 13175 10121 13201 10127
rect 13175 10089 13201 10095
rect 14855 10121 14881 10127
rect 14855 10089 14881 10095
rect 7687 10065 7713 10071
rect 7345 10039 7351 10065
rect 7377 10039 7383 10065
rect 7687 10033 7713 10039
rect 8807 10065 8833 10071
rect 12615 10065 12641 10071
rect 9361 10039 9367 10065
rect 9393 10039 9399 10065
rect 11657 10039 11663 10065
rect 11689 10039 11695 10065
rect 8807 10033 8833 10039
rect 12615 10033 12641 10039
rect 12783 10065 12809 10071
rect 12783 10033 12809 10039
rect 14071 10065 14097 10071
rect 14071 10033 14097 10039
rect 14127 10065 14153 10071
rect 14127 10033 14153 10039
rect 14351 10065 14377 10071
rect 14351 10033 14377 10039
rect 14407 10065 14433 10071
rect 14407 10033 14433 10039
rect 14967 10065 14993 10071
rect 14967 10033 14993 10039
rect 15247 10065 15273 10071
rect 15247 10033 15273 10039
rect 7183 10009 7209 10015
rect 7631 10009 7657 10015
rect 7513 9983 7519 10009
rect 7545 9983 7551 10009
rect 7183 9977 7209 9983
rect 7631 9977 7657 9983
rect 8919 10009 8945 10015
rect 13231 10009 13257 10015
rect 9473 9983 9479 10009
rect 9505 9983 9511 10009
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 8919 9977 8945 9983
rect 13231 9977 13257 9983
rect 13455 10009 13481 10015
rect 13455 9977 13481 9983
rect 13567 10009 13593 10015
rect 13567 9977 13593 9983
rect 13679 10009 13705 10015
rect 13679 9977 13705 9983
rect 13903 10009 13929 10015
rect 13903 9977 13929 9983
rect 13959 10009 13985 10015
rect 13959 9977 13985 9983
rect 14239 10009 14265 10015
rect 14239 9977 14265 9983
rect 15023 10009 15049 10015
rect 15023 9977 15049 9983
rect 15135 10009 15161 10015
rect 15135 9977 15161 9983
rect 15303 10009 15329 10015
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 15303 9977 15329 9983
rect 8975 9953 9001 9959
rect 13623 9953 13649 9959
rect 9417 9927 9423 9953
rect 9449 9927 9455 9953
rect 8975 9921 9001 9927
rect 13623 9921 13649 9927
rect 14631 9953 14657 9959
rect 14631 9921 14657 9927
rect 20007 9953 20033 9959
rect 20007 9921 20033 9927
rect 7905 9871 7911 9897
rect 7937 9871 7943 9897
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8863 9729 8889 9735
rect 8863 9697 8889 9703
rect 20007 9729 20033 9735
rect 20007 9697 20033 9703
rect 7127 9673 7153 9679
rect 9255 9673 9281 9679
rect 9081 9647 9087 9673
rect 9113 9647 9119 9673
rect 7127 9641 7153 9647
rect 9255 9641 9281 9647
rect 9591 9673 9617 9679
rect 9591 9641 9617 9647
rect 9983 9673 10009 9679
rect 13225 9647 13231 9673
rect 13257 9647 13263 9673
rect 14289 9647 14295 9673
rect 14321 9647 14327 9673
rect 9983 9641 10009 9647
rect 8135 9617 8161 9623
rect 8135 9585 8161 9591
rect 10039 9617 10065 9623
rect 10039 9585 10065 9591
rect 10207 9617 10233 9623
rect 10207 9585 10233 9591
rect 11159 9617 11185 9623
rect 11887 9617 11913 9623
rect 11433 9591 11439 9617
rect 11465 9591 11471 9617
rect 11159 9585 11185 9591
rect 11887 9585 11913 9591
rect 12167 9617 12193 9623
rect 12889 9591 12895 9617
rect 12921 9591 12927 9617
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 12167 9585 12193 9591
rect 8807 9561 8833 9567
rect 7569 9535 7575 9561
rect 7601 9535 7607 9561
rect 7905 9535 7911 9561
rect 7937 9535 7943 9561
rect 8807 9529 8833 9535
rect 9703 9561 9729 9567
rect 9703 9529 9729 9535
rect 9927 9561 9953 9567
rect 11271 9561 11297 9567
rect 10705 9535 10711 9561
rect 10737 9535 10743 9561
rect 10929 9535 10935 9561
rect 10961 9535 10967 9561
rect 9927 9529 9953 9535
rect 11271 9529 11297 9535
rect 12111 9561 12137 9567
rect 12111 9529 12137 9535
rect 7407 9505 7433 9511
rect 7407 9473 7433 9479
rect 7743 9505 7769 9511
rect 7743 9473 7769 9479
rect 8079 9505 8105 9511
rect 8079 9473 8105 9479
rect 8863 9505 8889 9511
rect 8863 9473 8889 9479
rect 9759 9505 9785 9511
rect 11775 9505 11801 9511
rect 11545 9479 11551 9505
rect 11577 9479 11583 9505
rect 9759 9473 9785 9479
rect 11775 9473 11801 9479
rect 11831 9505 11857 9511
rect 11831 9473 11857 9479
rect 11999 9505 12025 9511
rect 11999 9473 12025 9479
rect 14631 9505 14657 9511
rect 14631 9473 14657 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 10823 9337 10849 9343
rect 10823 9305 10849 9311
rect 12839 9337 12865 9343
rect 12839 9305 12865 9311
rect 9311 9281 9337 9287
rect 5945 9255 5951 9281
rect 5977 9255 5983 9281
rect 9311 9249 9337 9255
rect 9367 9281 9393 9287
rect 11489 9255 11495 9281
rect 11521 9255 11527 9281
rect 12945 9255 12951 9281
rect 12977 9255 12983 9281
rect 9367 9249 9393 9255
rect 7239 9225 7265 9231
rect 9871 9225 9897 9231
rect 10655 9225 10681 9231
rect 5609 9199 5615 9225
rect 5641 9199 5647 9225
rect 7401 9199 7407 9225
rect 7433 9199 7439 9225
rect 10145 9199 10151 9225
rect 10177 9199 10183 9225
rect 7239 9193 7265 9199
rect 9871 9193 9897 9199
rect 10655 9193 10681 9199
rect 10991 9225 11017 9231
rect 10991 9193 11017 9199
rect 11663 9225 11689 9231
rect 11663 9193 11689 9199
rect 12615 9225 12641 9231
rect 12615 9193 12641 9199
rect 13063 9225 13089 9231
rect 13399 9225 13425 9231
rect 13281 9199 13287 9225
rect 13313 9199 13319 9225
rect 13063 9193 13089 9199
rect 13399 9193 13425 9199
rect 13455 9225 13481 9231
rect 13455 9193 13481 9199
rect 7183 9169 7209 9175
rect 7009 9143 7015 9169
rect 7041 9143 7047 9169
rect 7183 9137 7209 9143
rect 9591 9169 9617 9175
rect 10201 9143 10207 9169
rect 10233 9143 10239 9169
rect 11209 9143 11215 9169
rect 11241 9143 11247 9169
rect 13113 9143 13119 9169
rect 13145 9143 13151 9169
rect 9591 9137 9617 9143
rect 9367 9113 9393 9119
rect 12671 9113 12697 9119
rect 10369 9087 10375 9113
rect 10401 9087 10407 9113
rect 13673 9087 13679 9113
rect 13705 9087 13711 9113
rect 9367 9081 9393 9087
rect 12671 9081 12697 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 12223 8945 12249 8951
rect 12223 8913 12249 8919
rect 14911 8945 14937 8951
rect 14911 8913 14937 8919
rect 12335 8889 12361 8895
rect 9193 8863 9199 8889
rect 9225 8863 9231 8889
rect 10257 8863 10263 8889
rect 10289 8863 10295 8889
rect 12335 8857 12361 8863
rect 12503 8889 12529 8895
rect 12503 8857 12529 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 7071 8833 7097 8839
rect 10711 8833 10737 8839
rect 8801 8807 8807 8833
rect 8833 8807 8839 8833
rect 7071 8801 7097 8807
rect 10711 8801 10737 8807
rect 11383 8833 11409 8839
rect 11383 8801 11409 8807
rect 11607 8833 11633 8839
rect 11607 8801 11633 8807
rect 12559 8833 12585 8839
rect 12895 8833 12921 8839
rect 12777 8807 12783 8833
rect 12809 8807 12815 8833
rect 12559 8801 12585 8807
rect 12895 8801 12921 8807
rect 12951 8833 12977 8839
rect 12951 8801 12977 8807
rect 13791 8833 13817 8839
rect 13791 8801 13817 8807
rect 14967 8833 14993 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 14967 8801 14993 8807
rect 6903 8777 6929 8783
rect 6903 8745 6929 8751
rect 11327 8777 11353 8783
rect 11327 8745 11353 8751
rect 11215 8721 11241 8727
rect 11215 8689 11241 8695
rect 11663 8721 11689 8727
rect 11663 8689 11689 8695
rect 11775 8721 11801 8727
rect 11775 8689 11801 8695
rect 12447 8721 12473 8727
rect 13959 8721 13985 8727
rect 13169 8695 13175 8721
rect 13201 8695 13207 8721
rect 12447 8689 12473 8695
rect 13959 8689 13985 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7295 8553 7321 8559
rect 7295 8521 7321 8527
rect 13399 8497 13425 8503
rect 6001 8471 6007 8497
rect 6033 8471 6039 8497
rect 9921 8471 9927 8497
rect 9953 8471 9959 8497
rect 13399 8465 13425 8471
rect 13567 8497 13593 8503
rect 14289 8471 14295 8497
rect 14321 8471 14327 8497
rect 13567 8465 13593 8471
rect 5609 8415 5615 8441
rect 5641 8415 5647 8441
rect 9809 8415 9815 8441
rect 9841 8415 9847 8441
rect 13897 8415 13903 8441
rect 13929 8415 13935 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 20007 8385 20033 8391
rect 7065 8359 7071 8385
rect 7097 8359 7103 8385
rect 15353 8359 15359 8385
rect 15385 8359 15391 8385
rect 20007 8353 20033 8359
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 11775 8161 11801 8167
rect 11775 8129 11801 8135
rect 14575 8161 14601 8167
rect 14575 8129 14601 8135
rect 8751 8105 8777 8111
rect 8751 8073 8777 8079
rect 8247 8049 8273 8055
rect 8247 8017 8273 8023
rect 8303 8049 8329 8055
rect 8975 8049 9001 8055
rect 8521 8023 8527 8049
rect 8553 8023 8559 8049
rect 8303 8017 8329 8023
rect 8975 8017 9001 8023
rect 9031 8049 9057 8055
rect 9031 8017 9057 8023
rect 9087 8049 9113 8055
rect 9087 8017 9113 8023
rect 11887 8049 11913 8055
rect 11993 8023 11999 8049
rect 12025 8023 12031 8049
rect 11887 8017 11913 8023
rect 12167 7993 12193 7999
rect 12167 7961 12193 7967
rect 14631 7993 14657 7999
rect 14631 7961 14657 7967
rect 8359 7937 8385 7943
rect 8359 7905 8385 7911
rect 8415 7937 8441 7943
rect 8415 7905 8441 7911
rect 8695 7937 8721 7943
rect 11943 7937 11969 7943
rect 9305 7911 9311 7937
rect 9337 7911 9343 7937
rect 8695 7905 8721 7911
rect 11943 7905 11969 7911
rect 12223 7937 12249 7943
rect 12223 7905 12249 7911
rect 12279 7937 12305 7943
rect 12279 7905 12305 7911
rect 13735 7937 13761 7943
rect 13735 7905 13761 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 9087 7769 9113 7775
rect 9087 7737 9113 7743
rect 12783 7769 12809 7775
rect 12783 7737 12809 7743
rect 15023 7769 15049 7775
rect 15023 7737 15049 7743
rect 8695 7713 8721 7719
rect 8695 7681 8721 7687
rect 8863 7713 8889 7719
rect 8863 7681 8889 7687
rect 9199 7713 9225 7719
rect 9199 7681 9225 7687
rect 9255 7713 9281 7719
rect 9255 7681 9281 7687
rect 10823 7713 10849 7719
rect 10823 7681 10849 7687
rect 10991 7713 11017 7719
rect 12945 7687 12951 7713
rect 12977 7687 12983 7713
rect 13729 7687 13735 7713
rect 13761 7687 13767 7713
rect 10991 7681 11017 7687
rect 8975 7657 9001 7663
rect 6897 7631 6903 7657
rect 6929 7631 6935 7657
rect 8975 7625 9001 7631
rect 11383 7657 11409 7663
rect 11383 7625 11409 7631
rect 11495 7657 11521 7663
rect 13337 7631 13343 7657
rect 13369 7631 13375 7657
rect 11495 7625 11521 7631
rect 8751 7601 8777 7607
rect 7233 7575 7239 7601
rect 7265 7575 7271 7601
rect 8297 7575 8303 7601
rect 8329 7575 8335 7601
rect 14793 7575 14799 7601
rect 14825 7575 14831 7601
rect 8751 7569 8777 7575
rect 11327 7545 11353 7551
rect 11327 7513 11353 7519
rect 11551 7545 11577 7551
rect 11551 7513 11577 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 8415 7377 8441 7383
rect 8415 7345 8441 7351
rect 9311 7377 9337 7383
rect 9311 7345 9337 7351
rect 9423 7377 9449 7383
rect 9423 7345 9449 7351
rect 9927 7377 9953 7383
rect 9927 7345 9953 7351
rect 10767 7377 10793 7383
rect 10767 7345 10793 7351
rect 10879 7377 10905 7383
rect 10879 7345 10905 7351
rect 11439 7377 11465 7383
rect 11439 7345 11465 7351
rect 8471 7321 8497 7327
rect 7177 7295 7183 7321
rect 7209 7295 7215 7321
rect 8241 7295 8247 7321
rect 8273 7295 8279 7321
rect 9753 7295 9759 7321
rect 9785 7295 9791 7321
rect 10369 7295 10375 7321
rect 10401 7295 10407 7321
rect 11993 7295 11999 7321
rect 12025 7295 12031 7321
rect 13057 7295 13063 7321
rect 13089 7295 13095 7321
rect 8471 7289 8497 7295
rect 8807 7265 8833 7271
rect 10207 7265 10233 7271
rect 11271 7265 11297 7271
rect 6841 7239 6847 7265
rect 6873 7239 6879 7265
rect 8577 7239 8583 7265
rect 8609 7239 8615 7265
rect 9529 7239 9535 7265
rect 9561 7239 9567 7265
rect 10649 7239 10655 7265
rect 10681 7239 10687 7265
rect 11433 7239 11439 7265
rect 11465 7239 11471 7265
rect 11601 7239 11607 7265
rect 11633 7239 11639 7265
rect 8807 7233 8833 7239
rect 10207 7233 10233 7239
rect 11271 7233 11297 7239
rect 9255 7209 9281 7215
rect 9255 7177 9281 7183
rect 9815 7153 9841 7159
rect 9815 7121 9841 7127
rect 10319 7153 10345 7159
rect 10319 7121 10345 7127
rect 10711 7153 10737 7159
rect 10711 7121 10737 7127
rect 13287 7153 13313 7159
rect 13287 7121 13313 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8359 6985 8385 6991
rect 8359 6953 8385 6959
rect 9641 6903 9647 6929
rect 9673 6903 9679 6929
rect 11265 6903 11271 6929
rect 11297 6903 11303 6929
rect 12671 6873 12697 6879
rect 9305 6847 9311 6873
rect 9337 6847 9343 6873
rect 10929 6847 10935 6873
rect 10961 6847 10967 6873
rect 12671 6841 12697 6847
rect 10705 6791 10711 6817
rect 10737 6791 10743 6817
rect 12329 6791 12335 6817
rect 12361 6791 12367 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 10319 6537 10345 6543
rect 8969 6511 8975 6537
rect 9001 6511 9007 6537
rect 10033 6511 10039 6537
rect 10065 6511 10071 6537
rect 10319 6505 10345 6511
rect 10823 6537 10849 6543
rect 10823 6505 10849 6511
rect 8577 6455 8583 6481
rect 8609 6455 8615 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 13399 2617 13425 2623
rect 13399 2585 13425 2591
rect 12889 2535 12895 2561
rect 12921 2535 12927 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8689 2143 8695 2169
rect 8721 2143 8727 2169
rect 10201 2143 10207 2169
rect 10233 2143 10239 2169
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 9249 2087 9255 2113
rect 9281 2087 9287 2113
rect 10711 2057 10737 2063
rect 10711 2025 10737 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 11215 1833 11241 1839
rect 11215 1801 11241 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8633 1751 8639 1777
rect 8665 1751 8671 1777
rect 10705 1751 10711 1777
rect 10737 1751 10743 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 9031 1665 9057 1671
rect 9031 1633 9057 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9031 19111 9057 19137
rect 11047 19111 11073 19137
rect 12783 19111 12809 19137
rect 14687 19111 14713 19137
rect 8527 18999 8553 19025
rect 10543 18999 10569 19025
rect 12279 18999 12305 19025
rect 14295 18999 14321 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10711 18719 10737 18745
rect 13399 18719 13425 18745
rect 10207 18607 10233 18633
rect 13119 18607 13145 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 967 13567 993 13593
rect 8527 13567 8553 13593
rect 10375 13567 10401 13593
rect 13175 13567 13201 13593
rect 20007 13567 20033 13593
rect 2143 13511 2169 13537
rect 7071 13511 7097 13537
rect 8919 13511 8945 13537
rect 11775 13511 11801 13537
rect 18943 13511 18969 13537
rect 7463 13455 7489 13481
rect 9311 13455 9337 13481
rect 12111 13455 12137 13481
rect 13399 13455 13425 13481
rect 8751 13399 8777 13425
rect 10711 13399 10737 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7855 13231 7881 13257
rect 12671 13231 12697 13257
rect 13119 13231 13145 13257
rect 8247 13175 8273 13201
rect 10431 13175 10457 13201
rect 12727 13175 12753 13201
rect 7463 13119 7489 13145
rect 7743 13119 7769 13145
rect 8023 13119 8049 13145
rect 8359 13119 8385 13145
rect 8751 13119 8777 13145
rect 10711 13119 10737 13145
rect 12335 13119 12361 13145
rect 12951 13119 12977 13145
rect 13455 13119 13481 13145
rect 18831 13119 18857 13145
rect 6063 13063 6089 13089
rect 7127 13063 7153 13089
rect 8135 13063 8161 13089
rect 9143 13063 9169 13089
rect 10207 13063 10233 13089
rect 11047 13063 11073 13089
rect 12111 13063 12137 13089
rect 13791 13063 13817 13089
rect 14855 13063 14881 13089
rect 15079 13063 15105 13089
rect 7911 13007 7937 13033
rect 12615 13007 12641 13033
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 7015 12839 7041 12865
rect 10263 12839 10289 12865
rect 11551 12839 11577 12865
rect 12615 12839 12641 12865
rect 13735 12839 13761 12865
rect 967 12783 993 12809
rect 10711 12783 10737 12809
rect 11271 12783 11297 12809
rect 2143 12727 2169 12753
rect 7855 12727 7881 12753
rect 9703 12727 9729 12753
rect 10039 12727 10065 12753
rect 10095 12727 10121 12753
rect 11103 12727 11129 12753
rect 11383 12727 11409 12753
rect 12335 12727 12361 12753
rect 14295 12727 14321 12753
rect 14799 12727 14825 12753
rect 6959 12671 6985 12697
rect 7519 12671 7545 12697
rect 7575 12671 7601 12697
rect 7631 12671 7657 12697
rect 9535 12671 9561 12697
rect 9983 12671 10009 12697
rect 10655 12671 10681 12697
rect 11159 12671 11185 12697
rect 11495 12671 11521 12697
rect 11551 12671 11577 12697
rect 12279 12671 12305 12697
rect 12391 12671 12417 12697
rect 12783 12671 12809 12697
rect 12839 12671 12865 12697
rect 12951 12671 12977 12697
rect 13791 12671 13817 12697
rect 14239 12671 14265 12697
rect 14519 12671 14545 12697
rect 14631 12671 14657 12697
rect 14687 12671 14713 12697
rect 14911 12671 14937 12697
rect 14967 12671 14993 12697
rect 7239 12615 7265 12641
rect 7463 12615 7489 12641
rect 8079 12615 8105 12641
rect 9591 12615 9617 12641
rect 9927 12615 9953 12641
rect 10767 12615 10793 12641
rect 13735 12615 13761 12641
rect 14127 12615 14153 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7351 12447 7377 12473
rect 9759 12447 9785 12473
rect 13679 12447 13705 12473
rect 6679 12391 6705 12417
rect 10263 12391 10289 12417
rect 14239 12391 14265 12417
rect 7071 12335 7097 12361
rect 7295 12335 7321 12361
rect 7407 12335 7433 12361
rect 7687 12335 7713 12361
rect 8639 12335 8665 12361
rect 8863 12335 8889 12361
rect 8975 12335 9001 12361
rect 9647 12335 9673 12361
rect 9983 12335 10009 12361
rect 10207 12335 10233 12361
rect 13847 12335 13873 12361
rect 18831 12335 18857 12361
rect 5615 12279 5641 12305
rect 8919 12279 8945 12305
rect 15303 12279 15329 12305
rect 7575 12223 7601 12249
rect 9815 12223 9841 12249
rect 10095 12223 10121 12249
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 7183 12055 7209 12081
rect 11103 12055 11129 12081
rect 7127 11999 7153 12025
rect 9535 11999 9561 12025
rect 10767 11999 10793 12025
rect 14295 11999 14321 12025
rect 16031 11999 16057 12025
rect 9255 11943 9281 11969
rect 9367 11943 9393 11969
rect 11047 11943 11073 11969
rect 11439 11943 11465 11969
rect 14575 11943 14601 11969
rect 8359 11887 8385 11913
rect 9815 11887 9841 11913
rect 9871 11887 9897 11913
rect 14967 11887 14993 11913
rect 7407 11831 7433 11857
rect 8527 11831 8553 11857
rect 9031 11831 9057 11857
rect 9983 11831 10009 11857
rect 10711 11831 10737 11857
rect 10823 11831 10849 11857
rect 11159 11831 11185 11857
rect 11271 11831 11297 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7799 11663 7825 11689
rect 8863 11663 8889 11689
rect 9367 11663 9393 11689
rect 10431 11663 10457 11689
rect 10655 11663 10681 11689
rect 11159 11663 11185 11689
rect 11775 11663 11801 11689
rect 12783 11663 12809 11689
rect 14687 11663 14713 11689
rect 14799 11663 14825 11689
rect 15191 11663 15217 11689
rect 8807 11607 8833 11633
rect 8975 11607 9001 11633
rect 9087 11607 9113 11633
rect 9535 11607 9561 11633
rect 9815 11607 9841 11633
rect 10319 11607 10345 11633
rect 10543 11607 10569 11633
rect 11831 11607 11857 11633
rect 13343 11607 13369 11633
rect 2143 11551 2169 11577
rect 7071 11551 7097 11577
rect 7351 11551 7377 11577
rect 7519 11551 7545 11577
rect 7631 11551 7657 11577
rect 7967 11551 7993 11577
rect 10263 11551 10289 11577
rect 10767 11551 10793 11577
rect 10991 11551 11017 11577
rect 11663 11551 11689 11577
rect 12671 11551 12697 11577
rect 13007 11551 13033 11577
rect 13231 11551 13257 11577
rect 13399 11551 13425 11577
rect 14855 11551 14881 11577
rect 15079 11551 15105 11577
rect 15247 11551 15273 11577
rect 5615 11495 5641 11521
rect 6679 11495 6705 11521
rect 7407 11495 7433 11521
rect 9759 11495 9785 11521
rect 10655 11495 10681 11521
rect 12727 11495 12753 11521
rect 967 11439 993 11465
rect 9703 11439 9729 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7183 11271 7209 11297
rect 9199 11215 9225 11241
rect 12727 11215 12753 11241
rect 13791 11215 13817 11241
rect 14015 11215 14041 11241
rect 20007 11215 20033 11241
rect 7239 11159 7265 11185
rect 7855 11159 7881 11185
rect 7911 11159 7937 11185
rect 9535 11159 9561 11185
rect 9703 11159 9729 11185
rect 10767 11159 10793 11185
rect 11047 11159 11073 11185
rect 11103 11159 11129 11185
rect 11327 11159 11353 11185
rect 11999 11159 12025 11185
rect 12391 11159 12417 11185
rect 18831 11159 18857 11185
rect 7183 11103 7209 11129
rect 7631 11103 7657 11129
rect 7743 11103 7769 11129
rect 9479 11103 9505 11129
rect 9983 11103 10009 11129
rect 10991 11103 11017 11129
rect 11495 11103 11521 11129
rect 12055 11103 12081 11129
rect 7687 11047 7713 11073
rect 10655 11047 10681 11073
rect 12167 11047 12193 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8415 10879 8441 10905
rect 11943 10879 11969 10905
rect 14911 10879 14937 10905
rect 6063 10823 6089 10849
rect 9255 10823 9281 10849
rect 11551 10823 11577 10849
rect 14687 10823 14713 10849
rect 5671 10767 5697 10793
rect 8303 10767 8329 10793
rect 11327 10767 11353 10793
rect 11495 10767 11521 10793
rect 11663 10767 11689 10793
rect 12111 10767 12137 10793
rect 12895 10767 12921 10793
rect 14519 10767 14545 10793
rect 18831 10767 18857 10793
rect 7127 10711 7153 10737
rect 7351 10711 7377 10737
rect 13287 10711 13313 10737
rect 14351 10711 14377 10737
rect 20007 10711 20033 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7519 10487 7545 10513
rect 10039 10487 10065 10513
rect 10319 10487 10345 10513
rect 10655 10487 10681 10513
rect 7967 10431 7993 10457
rect 9479 10431 9505 10457
rect 10935 10431 10961 10457
rect 12895 10431 12921 10457
rect 16087 10431 16113 10457
rect 20007 10431 20033 10457
rect 7463 10375 7489 10401
rect 8247 10375 8273 10401
rect 8527 10375 8553 10401
rect 8639 10375 8665 10401
rect 8807 10375 8833 10401
rect 9255 10375 9281 10401
rect 9759 10375 9785 10401
rect 10375 10375 10401 10401
rect 10823 10375 10849 10401
rect 11103 10375 11129 10401
rect 11215 10375 11241 10401
rect 11663 10375 11689 10401
rect 14631 10375 14657 10401
rect 16311 10375 16337 10401
rect 18831 10375 18857 10401
rect 8359 10319 8385 10345
rect 9983 10319 10009 10345
rect 10151 10319 10177 10345
rect 15023 10319 15049 10345
rect 16423 10319 16449 10345
rect 7687 10263 7713 10289
rect 8583 10263 8609 10289
rect 9871 10263 9897 10289
rect 10263 10263 10289 10289
rect 11159 10263 11185 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 8079 10095 8105 10121
rect 8247 10095 8273 10121
rect 9031 10095 9057 10121
rect 13119 10095 13145 10121
rect 13175 10095 13201 10121
rect 14855 10095 14881 10121
rect 7351 10039 7377 10065
rect 7687 10039 7713 10065
rect 8807 10039 8833 10065
rect 9367 10039 9393 10065
rect 11663 10039 11689 10065
rect 12615 10039 12641 10065
rect 12783 10039 12809 10065
rect 14071 10039 14097 10065
rect 14127 10039 14153 10065
rect 14351 10039 14377 10065
rect 14407 10039 14433 10065
rect 14967 10039 14993 10065
rect 15247 10039 15273 10065
rect 7183 9983 7209 10009
rect 7519 9983 7545 10009
rect 7631 9983 7657 10009
rect 8919 9983 8945 10009
rect 9479 9983 9505 10009
rect 9703 9983 9729 10009
rect 13231 9983 13257 10009
rect 13455 9983 13481 10009
rect 13567 9983 13593 10009
rect 13679 9983 13705 10009
rect 13903 9983 13929 10009
rect 13959 9983 13985 10009
rect 14239 9983 14265 10009
rect 15023 9983 15049 10009
rect 15135 9983 15161 10009
rect 15303 9983 15329 10009
rect 18831 9983 18857 10009
rect 8975 9927 9001 9953
rect 9423 9927 9449 9953
rect 13623 9927 13649 9953
rect 14631 9927 14657 9953
rect 20007 9927 20033 9953
rect 7911 9871 7937 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8863 9703 8889 9729
rect 20007 9703 20033 9729
rect 7127 9647 7153 9673
rect 9087 9647 9113 9673
rect 9255 9647 9281 9673
rect 9591 9647 9617 9673
rect 9983 9647 10009 9673
rect 13231 9647 13257 9673
rect 14295 9647 14321 9673
rect 8135 9591 8161 9617
rect 10039 9591 10065 9617
rect 10207 9591 10233 9617
rect 11159 9591 11185 9617
rect 11439 9591 11465 9617
rect 11887 9591 11913 9617
rect 12167 9591 12193 9617
rect 12895 9591 12921 9617
rect 18831 9591 18857 9617
rect 7575 9535 7601 9561
rect 7911 9535 7937 9561
rect 8807 9535 8833 9561
rect 9703 9535 9729 9561
rect 9927 9535 9953 9561
rect 10711 9535 10737 9561
rect 10935 9535 10961 9561
rect 11271 9535 11297 9561
rect 12111 9535 12137 9561
rect 7407 9479 7433 9505
rect 7743 9479 7769 9505
rect 8079 9479 8105 9505
rect 8863 9479 8889 9505
rect 9759 9479 9785 9505
rect 11551 9479 11577 9505
rect 11775 9479 11801 9505
rect 11831 9479 11857 9505
rect 11999 9479 12025 9505
rect 14631 9479 14657 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 10823 9311 10849 9337
rect 12839 9311 12865 9337
rect 5951 9255 5977 9281
rect 9311 9255 9337 9281
rect 9367 9255 9393 9281
rect 11495 9255 11521 9281
rect 12951 9255 12977 9281
rect 5615 9199 5641 9225
rect 7239 9199 7265 9225
rect 7407 9199 7433 9225
rect 9871 9199 9897 9225
rect 10151 9199 10177 9225
rect 10655 9199 10681 9225
rect 10991 9199 11017 9225
rect 11663 9199 11689 9225
rect 12615 9199 12641 9225
rect 13063 9199 13089 9225
rect 13287 9199 13313 9225
rect 13399 9199 13425 9225
rect 13455 9199 13481 9225
rect 7015 9143 7041 9169
rect 7183 9143 7209 9169
rect 9591 9143 9617 9169
rect 10207 9143 10233 9169
rect 11215 9143 11241 9169
rect 13119 9143 13145 9169
rect 9367 9087 9393 9113
rect 10375 9087 10401 9113
rect 12671 9087 12697 9113
rect 13679 9087 13705 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 12223 8919 12249 8945
rect 14911 8919 14937 8945
rect 9199 8863 9225 8889
rect 10263 8863 10289 8889
rect 12335 8863 12361 8889
rect 12503 8863 12529 8889
rect 20007 8863 20033 8889
rect 7071 8807 7097 8833
rect 8807 8807 8833 8833
rect 10711 8807 10737 8833
rect 11383 8807 11409 8833
rect 11607 8807 11633 8833
rect 12559 8807 12585 8833
rect 12783 8807 12809 8833
rect 12895 8807 12921 8833
rect 12951 8807 12977 8833
rect 13791 8807 13817 8833
rect 14967 8807 14993 8833
rect 18831 8807 18857 8833
rect 6903 8751 6929 8777
rect 11327 8751 11353 8777
rect 11215 8695 11241 8721
rect 11663 8695 11689 8721
rect 11775 8695 11801 8721
rect 12447 8695 12473 8721
rect 13175 8695 13201 8721
rect 13959 8695 13985 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7295 8527 7321 8553
rect 6007 8471 6033 8497
rect 9927 8471 9953 8497
rect 13399 8471 13425 8497
rect 13567 8471 13593 8497
rect 14295 8471 14321 8497
rect 5615 8415 5641 8441
rect 9815 8415 9841 8441
rect 13903 8415 13929 8441
rect 18831 8415 18857 8441
rect 7071 8359 7097 8385
rect 15359 8359 15385 8385
rect 20007 8359 20033 8385
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 11775 8135 11801 8161
rect 14575 8135 14601 8161
rect 8751 8079 8777 8105
rect 8247 8023 8273 8049
rect 8303 8023 8329 8049
rect 8527 8023 8553 8049
rect 8975 8023 9001 8049
rect 9031 8023 9057 8049
rect 9087 8023 9113 8049
rect 11887 8023 11913 8049
rect 11999 8023 12025 8049
rect 12167 7967 12193 7993
rect 14631 7967 14657 7993
rect 8359 7911 8385 7937
rect 8415 7911 8441 7937
rect 8695 7911 8721 7937
rect 9311 7911 9337 7937
rect 11943 7911 11969 7937
rect 12223 7911 12249 7937
rect 12279 7911 12305 7937
rect 13735 7911 13761 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 9087 7743 9113 7769
rect 12783 7743 12809 7769
rect 15023 7743 15049 7769
rect 8695 7687 8721 7713
rect 8863 7687 8889 7713
rect 9199 7687 9225 7713
rect 9255 7687 9281 7713
rect 10823 7687 10849 7713
rect 10991 7687 11017 7713
rect 12951 7687 12977 7713
rect 13735 7687 13761 7713
rect 6903 7631 6929 7657
rect 8975 7631 9001 7657
rect 11383 7631 11409 7657
rect 11495 7631 11521 7657
rect 13343 7631 13369 7657
rect 7239 7575 7265 7601
rect 8303 7575 8329 7601
rect 8751 7575 8777 7601
rect 14799 7575 14825 7601
rect 11327 7519 11353 7545
rect 11551 7519 11577 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8415 7351 8441 7377
rect 9311 7351 9337 7377
rect 9423 7351 9449 7377
rect 9927 7351 9953 7377
rect 10767 7351 10793 7377
rect 10879 7351 10905 7377
rect 11439 7351 11465 7377
rect 7183 7295 7209 7321
rect 8247 7295 8273 7321
rect 8471 7295 8497 7321
rect 9759 7295 9785 7321
rect 10375 7295 10401 7321
rect 11999 7295 12025 7321
rect 13063 7295 13089 7321
rect 6847 7239 6873 7265
rect 8583 7239 8609 7265
rect 8807 7239 8833 7265
rect 9535 7239 9561 7265
rect 10207 7239 10233 7265
rect 10655 7239 10681 7265
rect 11271 7239 11297 7265
rect 11439 7239 11465 7265
rect 11607 7239 11633 7265
rect 9255 7183 9281 7209
rect 9815 7127 9841 7153
rect 10319 7127 10345 7153
rect 10711 7127 10737 7153
rect 13287 7127 13313 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8359 6959 8385 6985
rect 9647 6903 9673 6929
rect 11271 6903 11297 6929
rect 9311 6847 9337 6873
rect 10935 6847 10961 6873
rect 12671 6847 12697 6873
rect 10711 6791 10737 6817
rect 12335 6791 12361 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8975 6511 9001 6537
rect 10039 6511 10065 6537
rect 10319 6511 10345 6537
rect 10823 6511 10849 6537
rect 8583 6455 8609 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 13399 2591 13425 2617
rect 12895 2535 12921 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8695 2143 8721 2169
rect 10207 2143 10233 2169
rect 12615 2143 12641 2169
rect 9255 2087 9281 2113
rect 10711 2031 10737 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 11215 1807 11241 1833
rect 12783 1807 12809 1833
rect 8639 1751 8665 1777
rect 10711 1751 10737 1777
rect 12279 1751 12305 1777
rect 9031 1639 9057 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 12096 20600 12152 21000
rect 12768 20600 12824 21000
rect 13104 20600 13160 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8414 19138 8442 20600
rect 8414 19105 8442 19110
rect 9030 19138 9058 19143
rect 9030 19091 9058 19110
rect 8526 19025 8554 19031
rect 8526 18999 8527 19025
rect 8553 18999 8554 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 966 13593 994 13599
rect 8526 13594 8554 18999
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10094 18746 10122 20600
rect 10430 19138 10458 20600
rect 10430 19105 10458 19110
rect 11046 19138 11074 19143
rect 11046 19091 11074 19110
rect 12110 19138 12138 20600
rect 12782 19306 12810 20600
rect 12782 19273 12810 19278
rect 12110 19105 12138 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 13118 19138 13146 20600
rect 13118 19105 13146 19110
rect 13398 19306 13426 19311
rect 10094 18713 10122 18718
rect 10542 19025 10570 19031
rect 10542 18999 10543 19025
rect 10569 18999 10570 19025
rect 10206 18633 10234 18639
rect 10206 18607 10207 18633
rect 10233 18607 10234 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 966 13567 967 13593
rect 993 13567 994 13593
rect 966 13146 994 13567
rect 8414 13593 8554 13594
rect 8414 13567 8527 13593
rect 8553 13567 8554 13593
rect 8414 13566 8554 13567
rect 2142 13538 2170 13543
rect 2142 13491 2170 13510
rect 6062 13538 6090 13543
rect 966 13113 994 13118
rect 2086 13482 2114 13487
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 2086 9506 2114 13454
rect 6062 13090 6090 13510
rect 7070 13537 7098 13543
rect 7070 13511 7071 13537
rect 7097 13511 7098 13537
rect 7070 13202 7098 13511
rect 7462 13481 7490 13487
rect 7462 13455 7463 13481
rect 7489 13455 7490 13481
rect 7462 13426 7490 13455
rect 8414 13454 8442 13566
rect 8526 13561 8554 13566
rect 7462 13393 7490 13398
rect 7854 13426 7882 13431
rect 7854 13257 7882 13398
rect 7854 13231 7855 13257
rect 7881 13231 7882 13257
rect 7854 13225 7882 13231
rect 8246 13426 8442 13454
rect 8918 13537 8946 13543
rect 8918 13511 8919 13537
rect 8945 13511 8946 13537
rect 8750 13426 8778 13431
rect 8918 13426 8946 13511
rect 7070 13169 7098 13174
rect 7406 13202 7434 13207
rect 7406 13146 7434 13174
rect 8246 13201 8274 13426
rect 8246 13175 8247 13201
rect 8273 13175 8274 13201
rect 8246 13169 8274 13175
rect 8750 13425 8946 13426
rect 8750 13399 8751 13425
rect 8777 13399 8946 13425
rect 8750 13398 8946 13399
rect 9310 13481 9338 13487
rect 9310 13455 9311 13481
rect 9337 13455 9338 13481
rect 8750 13202 8778 13398
rect 7462 13146 7490 13151
rect 7742 13146 7770 13151
rect 8022 13146 8050 13151
rect 7406 13145 7490 13146
rect 7406 13119 7463 13145
rect 7489 13119 7490 13145
rect 7406 13118 7490 13119
rect 7126 13090 7154 13095
rect 6062 13043 6090 13062
rect 7014 13089 7154 13090
rect 7014 13063 7127 13089
rect 7153 13063 7154 13089
rect 7014 13062 7154 13063
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 7014 12865 7042 13062
rect 7126 13057 7154 13062
rect 7014 12839 7015 12865
rect 7041 12839 7042 12865
rect 7014 12833 7042 12839
rect 2142 12753 2170 12759
rect 2142 12727 2143 12753
rect 2169 12727 2170 12753
rect 2142 12306 2170 12727
rect 6958 12698 6986 12703
rect 6958 12651 6986 12670
rect 7238 12642 7266 12647
rect 7406 12642 7434 13118
rect 7462 13113 7490 13118
rect 7686 13145 7770 13146
rect 7686 13119 7743 13145
rect 7769 13119 7770 13145
rect 7686 13118 7770 13119
rect 7574 13090 7602 13095
rect 7518 12698 7546 12703
rect 7518 12651 7546 12670
rect 7574 12697 7602 13062
rect 7574 12671 7575 12697
rect 7601 12671 7602 12697
rect 7574 12665 7602 12671
rect 7630 12698 7658 12703
rect 7630 12651 7658 12670
rect 7238 12641 7406 12642
rect 7238 12615 7239 12641
rect 7265 12615 7406 12641
rect 7238 12614 7406 12615
rect 6678 12474 6706 12479
rect 6678 12417 6706 12446
rect 6678 12391 6679 12417
rect 6705 12391 6706 12417
rect 6678 12385 6706 12391
rect 7070 12362 7098 12367
rect 7238 12362 7266 12614
rect 7406 12595 7434 12614
rect 7462 12641 7490 12647
rect 7462 12615 7463 12641
rect 7489 12615 7490 12641
rect 7462 12586 7490 12615
rect 7686 12586 7714 13118
rect 7742 13113 7770 13118
rect 7854 13145 8050 13146
rect 7854 13119 8023 13145
rect 8049 13119 8050 13145
rect 7854 13118 8050 13119
rect 7462 12558 7686 12586
rect 7350 12474 7378 12479
rect 7350 12427 7378 12446
rect 7070 12361 7266 12362
rect 7070 12335 7071 12361
rect 7097 12335 7266 12361
rect 7070 12334 7266 12335
rect 7294 12362 7322 12367
rect 7406 12362 7434 12367
rect 2142 12273 2170 12278
rect 5614 12306 5642 12311
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 5614 12026 5642 12278
rect 5614 11993 5642 11998
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 7070 11578 7098 12334
rect 7294 12315 7322 12334
rect 7350 12361 7434 12362
rect 7350 12335 7407 12361
rect 7433 12335 7434 12361
rect 7350 12334 7434 12335
rect 7182 12082 7210 12087
rect 7350 12082 7378 12334
rect 7406 12329 7434 12334
rect 7574 12249 7602 12558
rect 7686 12539 7714 12558
rect 7854 12753 7882 13118
rect 8022 13113 8050 13118
rect 8358 13145 8386 13151
rect 8358 13119 8359 13145
rect 8385 13119 8386 13145
rect 8134 13089 8162 13095
rect 8134 13063 8135 13089
rect 8161 13063 8162 13089
rect 7910 13034 7938 13039
rect 8134 13034 8162 13063
rect 7910 13033 8162 13034
rect 7910 13007 7911 13033
rect 7937 13007 8162 13033
rect 7910 13006 8162 13007
rect 7910 13001 7938 13006
rect 7854 12727 7855 12753
rect 7881 12727 7882 12753
rect 7854 12474 7882 12727
rect 8078 12642 8106 12647
rect 8078 12595 8106 12614
rect 7574 12223 7575 12249
rect 7601 12223 7602 12249
rect 7574 12217 7602 12223
rect 7686 12361 7714 12367
rect 7686 12335 7687 12361
rect 7713 12335 7714 12361
rect 7182 12081 7378 12082
rect 7182 12055 7183 12081
rect 7209 12055 7378 12081
rect 7182 12054 7378 12055
rect 7182 12049 7210 12054
rect 7126 12026 7154 12031
rect 7126 11979 7154 11998
rect 7406 11858 7434 11863
rect 7294 11857 7434 11858
rect 7294 11831 7407 11857
rect 7433 11831 7434 11857
rect 7294 11830 7434 11831
rect 7294 11578 7322 11830
rect 7406 11825 7434 11830
rect 7686 11690 7714 12335
rect 7686 11657 7714 11662
rect 7798 11690 7826 11695
rect 7854 11690 7882 12446
rect 8302 12586 8330 12591
rect 8358 12586 8386 13119
rect 8750 13145 8778 13174
rect 8750 13119 8751 13145
rect 8777 13119 8778 13145
rect 8750 12642 8778 13119
rect 8750 12609 8778 12614
rect 9142 13089 9170 13095
rect 9142 13063 9143 13089
rect 9169 13063 9170 13089
rect 8638 12586 8666 12591
rect 8358 12558 8442 12586
rect 8022 12362 8050 12367
rect 7798 11689 7882 11690
rect 7798 11663 7799 11689
rect 7825 11663 7882 11689
rect 7798 11662 7882 11663
rect 7910 11690 7938 11695
rect 7070 11577 7322 11578
rect 7070 11551 7071 11577
rect 7097 11551 7322 11577
rect 7070 11550 7322 11551
rect 7350 11577 7378 11583
rect 7350 11551 7351 11577
rect 7377 11551 7378 11577
rect 5614 11522 5642 11527
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 5614 11130 5642 11494
rect 6678 11522 6706 11527
rect 6678 11475 6706 11494
rect 5614 11097 5642 11102
rect 6062 11074 6090 11079
rect 6062 10849 6090 11046
rect 7070 11018 7098 11550
rect 7350 11354 7378 11551
rect 7518 11577 7546 11583
rect 7518 11551 7519 11577
rect 7545 11551 7546 11577
rect 7406 11522 7434 11527
rect 7406 11475 7434 11494
rect 7182 11326 7378 11354
rect 7182 11297 7210 11326
rect 7182 11271 7183 11297
rect 7209 11271 7210 11297
rect 7182 11265 7210 11271
rect 7238 11186 7266 11191
rect 7238 11139 7266 11158
rect 7182 11130 7210 11135
rect 7518 11130 7546 11551
rect 7630 11577 7658 11583
rect 7630 11551 7631 11577
rect 7657 11551 7658 11577
rect 7630 11298 7658 11551
rect 7630 11265 7658 11270
rect 7798 11186 7826 11662
rect 7798 11153 7826 11158
rect 7854 11242 7882 11247
rect 7854 11185 7882 11214
rect 7854 11159 7855 11185
rect 7881 11159 7882 11185
rect 7630 11130 7658 11135
rect 7518 11129 7658 11130
rect 7518 11103 7631 11129
rect 7657 11103 7658 11129
rect 7518 11102 7658 11103
rect 7182 11083 7210 11102
rect 7070 10990 7210 11018
rect 6062 10823 6063 10849
rect 6089 10823 6090 10849
rect 6062 10817 6090 10823
rect 5670 10793 5698 10799
rect 5670 10767 5671 10793
rect 5697 10767 5698 10793
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 5670 10122 5698 10767
rect 7126 10738 7154 10743
rect 7182 10738 7210 10990
rect 7350 10850 7378 10855
rect 7350 10738 7378 10822
rect 7182 10737 7378 10738
rect 7182 10711 7351 10737
rect 7377 10711 7378 10737
rect 7182 10710 7378 10711
rect 7126 10691 7154 10710
rect 5614 10066 5698 10094
rect 7238 10122 7266 10127
rect 7294 10122 7322 10710
rect 7350 10705 7378 10710
rect 7462 10738 7490 10743
rect 7462 10402 7490 10710
rect 7518 10514 7546 10519
rect 7518 10467 7546 10486
rect 7630 10402 7658 11102
rect 7742 11129 7770 11135
rect 7742 11103 7743 11129
rect 7769 11103 7770 11129
rect 7686 11074 7714 11079
rect 7686 11027 7714 11046
rect 7742 10514 7770 11103
rect 7742 10481 7770 10486
rect 7462 10401 7602 10402
rect 7462 10375 7463 10401
rect 7489 10375 7602 10401
rect 7462 10374 7602 10375
rect 7630 10374 7770 10402
rect 7462 10369 7490 10374
rect 7574 10290 7602 10374
rect 7686 10290 7714 10295
rect 7574 10289 7714 10290
rect 7574 10263 7687 10289
rect 7713 10263 7714 10289
rect 7574 10262 7714 10263
rect 7266 10094 7322 10122
rect 7686 10122 7714 10262
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 2086 9473 2114 9478
rect 5614 9225 5642 10066
rect 7182 10010 7210 10015
rect 7014 10009 7210 10010
rect 7014 9983 7183 10009
rect 7209 9983 7210 10009
rect 7014 9982 7210 9983
rect 5950 9282 5978 9287
rect 5950 9235 5978 9254
rect 5614 9199 5615 9225
rect 5641 9199 5642 9225
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 5614 8441 5642 9199
rect 7014 9170 7042 9982
rect 7182 9977 7210 9982
rect 7126 9674 7154 9679
rect 7238 9674 7266 10094
rect 7350 10066 7378 10071
rect 7350 10019 7378 10038
rect 7686 10065 7714 10094
rect 7686 10039 7687 10065
rect 7713 10039 7714 10065
rect 7686 10033 7714 10039
rect 7518 10009 7546 10015
rect 7518 9983 7519 10009
rect 7545 9983 7546 10009
rect 7126 9673 7322 9674
rect 7126 9647 7127 9673
rect 7153 9647 7322 9673
rect 7126 9646 7322 9647
rect 7126 9641 7154 9646
rect 7238 9338 7266 9343
rect 7238 9225 7266 9310
rect 7238 9199 7239 9225
rect 7265 9199 7266 9225
rect 7182 9170 7210 9175
rect 7014 9123 7042 9142
rect 7070 9169 7210 9170
rect 7070 9143 7183 9169
rect 7209 9143 7210 9169
rect 7070 9142 7210 9143
rect 7070 8833 7098 9142
rect 7182 9137 7210 9142
rect 7070 8807 7071 8833
rect 7097 8807 7098 8833
rect 7070 8801 7098 8807
rect 6006 8778 6034 8783
rect 6006 8497 6034 8750
rect 6902 8778 6930 8783
rect 6902 8731 6930 8750
rect 6006 8471 6007 8497
rect 6033 8471 6034 8497
rect 6006 8465 6034 8471
rect 5614 8415 5615 8441
rect 5641 8415 5642 8441
rect 5614 8409 5642 8415
rect 7070 8386 7098 8391
rect 7238 8386 7266 9199
rect 7070 8385 7266 8386
rect 7070 8359 7071 8385
rect 7097 8359 7266 8385
rect 7070 8358 7266 8359
rect 7294 8553 7322 9646
rect 7406 9505 7434 9511
rect 7406 9479 7407 9505
rect 7433 9479 7434 9505
rect 7406 9338 7434 9479
rect 7406 9305 7434 9310
rect 7406 9226 7434 9231
rect 7518 9226 7546 9983
rect 7630 10010 7658 10015
rect 7574 9562 7602 9567
rect 7630 9562 7658 9982
rect 7742 9898 7770 10374
rect 7854 9898 7882 11159
rect 7910 11185 7938 11662
rect 7910 11159 7911 11185
rect 7937 11159 7938 11185
rect 7910 11153 7938 11159
rect 7966 11577 7994 11583
rect 7966 11551 7967 11577
rect 7993 11551 7994 11577
rect 7966 11186 7994 11551
rect 8022 11242 8050 12334
rect 8302 11914 8330 12558
rect 8414 12530 8442 12558
rect 8470 12530 8498 12535
rect 8414 12502 8470 12530
rect 8470 12497 8498 12502
rect 8638 12361 8666 12558
rect 9030 12530 9058 12535
rect 8638 12335 8639 12361
rect 8665 12335 8666 12361
rect 8638 12329 8666 12335
rect 8862 12362 8890 12367
rect 8862 12315 8890 12334
rect 8974 12362 9002 12367
rect 9030 12362 9058 12502
rect 9142 12474 9170 13063
rect 9310 12866 9338 13455
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9310 12833 9338 12838
rect 10206 13089 10234 18607
rect 10542 15974 10570 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 10710 18746 10738 18751
rect 10710 18699 10738 18718
rect 12278 15974 12306 18999
rect 13398 18745 13426 19278
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 14686 19138 14714 19143
rect 14686 19091 14714 19110
rect 13398 18719 13399 18745
rect 13425 18719 13426 18745
rect 13398 18713 13426 18719
rect 14294 19025 14322 19031
rect 14294 18999 14295 19025
rect 14321 18999 14322 19025
rect 13118 18634 13146 18639
rect 13118 18633 13202 18634
rect 13118 18607 13119 18633
rect 13145 18607 13202 18633
rect 13118 18606 13202 18607
rect 13118 18601 13146 18606
rect 10374 15946 10570 15974
rect 12054 15946 12306 15974
rect 10374 13594 10402 15946
rect 10206 13063 10207 13089
rect 10233 13063 10234 13089
rect 10150 12810 10178 12815
rect 9814 12782 10066 12810
rect 9702 12754 9730 12759
rect 9702 12707 9730 12726
rect 9142 12441 9170 12446
rect 9198 12698 9226 12703
rect 8974 12361 9058 12362
rect 8974 12335 8975 12361
rect 9001 12335 9058 12361
rect 8974 12334 9058 12335
rect 8974 12329 9002 12334
rect 8918 12305 8946 12311
rect 8918 12279 8919 12305
rect 8945 12279 8946 12305
rect 8806 11970 8834 11975
rect 8358 11914 8386 11919
rect 8302 11913 8386 11914
rect 8302 11887 8359 11913
rect 8385 11887 8386 11913
rect 8302 11886 8386 11887
rect 8358 11881 8386 11886
rect 8526 11858 8554 11863
rect 8526 11811 8554 11830
rect 8806 11634 8834 11942
rect 8918 11746 8946 12279
rect 9030 11857 9058 12334
rect 9030 11831 9031 11857
rect 9057 11831 9058 11857
rect 9030 11825 9058 11831
rect 9086 11914 9114 11919
rect 8918 11713 8946 11718
rect 8862 11690 8890 11695
rect 8862 11643 8890 11662
rect 8022 11209 8050 11214
rect 8414 11633 8834 11634
rect 8414 11607 8807 11633
rect 8833 11607 8834 11633
rect 8414 11606 8834 11607
rect 7966 11130 7994 11158
rect 7966 11102 8050 11130
rect 7966 10458 7994 10463
rect 8022 10458 8050 11102
rect 8358 10906 8386 10911
rect 8302 10878 8358 10906
rect 8302 10793 8330 10878
rect 8358 10873 8386 10878
rect 8414 10905 8442 11606
rect 8414 10879 8415 10905
rect 8441 10879 8442 10905
rect 8414 10873 8442 10879
rect 8302 10767 8303 10793
rect 8329 10767 8330 10793
rect 7966 10457 8050 10458
rect 7966 10431 7967 10457
rect 7993 10431 8050 10457
rect 7966 10430 8050 10431
rect 8134 10570 8162 10575
rect 7966 10425 7994 10430
rect 8078 10122 8106 10127
rect 8078 10075 8106 10094
rect 8134 10066 8162 10542
rect 7910 9898 7938 9903
rect 7854 9897 7938 9898
rect 7854 9871 7911 9897
rect 7937 9871 7938 9897
rect 7854 9870 7938 9871
rect 7742 9865 7770 9870
rect 7910 9674 7938 9870
rect 7910 9641 7938 9646
rect 8134 9617 8162 10038
rect 8246 10401 8274 10407
rect 8246 10375 8247 10401
rect 8273 10375 8274 10401
rect 8246 10121 8274 10375
rect 8246 10095 8247 10121
rect 8273 10095 8274 10121
rect 8246 10066 8274 10095
rect 8246 10033 8274 10038
rect 8302 10010 8330 10767
rect 8750 10850 8778 10855
rect 8526 10402 8554 10407
rect 8358 10374 8526 10402
rect 8358 10345 8386 10374
rect 8526 10355 8554 10374
rect 8638 10401 8666 10407
rect 8638 10375 8639 10401
rect 8665 10375 8666 10401
rect 8358 10319 8359 10345
rect 8385 10319 8386 10345
rect 8358 10313 8386 10319
rect 8302 9977 8330 9982
rect 8582 10289 8610 10295
rect 8582 10263 8583 10289
rect 8609 10263 8610 10289
rect 8134 9591 8135 9617
rect 8161 9591 8162 9617
rect 8134 9585 8162 9591
rect 7574 9561 7658 9562
rect 7574 9535 7575 9561
rect 7601 9535 7658 9561
rect 7574 9534 7658 9535
rect 7910 9562 7938 9567
rect 7574 9529 7602 9534
rect 7910 9515 7938 9534
rect 7742 9505 7770 9511
rect 7742 9479 7743 9505
rect 7769 9479 7770 9505
rect 7742 9338 7770 9479
rect 7742 9305 7770 9310
rect 8078 9505 8106 9511
rect 8078 9479 8079 9505
rect 8105 9479 8106 9505
rect 8078 9282 8106 9479
rect 8078 9249 8106 9254
rect 7406 9225 7546 9226
rect 7406 9199 7407 9225
rect 7433 9199 7546 9225
rect 7406 9198 7546 9199
rect 7350 9170 7378 9175
rect 7406 9170 7434 9198
rect 7378 9142 7434 9170
rect 8246 9170 8274 9175
rect 7350 9137 7378 9142
rect 7294 8527 7295 8553
rect 7321 8527 7322 8553
rect 7070 8353 7098 8358
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 7294 7714 7322 8527
rect 8246 8049 8274 9142
rect 8582 9114 8610 10263
rect 8638 10010 8666 10375
rect 8638 9977 8666 9982
rect 8246 8023 8247 8049
rect 8273 8023 8274 8049
rect 8246 8017 8274 8023
rect 8302 9086 8610 9114
rect 8302 8049 8330 9086
rect 8750 8834 8778 10822
rect 8806 10401 8834 11606
rect 8974 11634 9002 11639
rect 8974 11587 9002 11606
rect 9086 11633 9114 11886
rect 9086 11607 9087 11633
rect 9113 11607 9114 11633
rect 8806 10375 8807 10401
rect 8833 10375 8834 10401
rect 8806 10369 8834 10375
rect 9030 11242 9058 11247
rect 9030 10122 9058 11214
rect 9086 10402 9114 11607
rect 9086 10369 9114 10374
rect 9198 11241 9226 12670
rect 9534 12697 9562 12703
rect 9534 12671 9535 12697
rect 9561 12671 9562 12697
rect 9534 12530 9562 12671
rect 9534 12497 9562 12502
rect 9590 12641 9618 12647
rect 9590 12615 9591 12641
rect 9617 12615 9618 12641
rect 9590 12474 9618 12615
rect 9758 12642 9786 12647
rect 9590 12446 9730 12474
rect 9254 12418 9282 12423
rect 9254 11970 9282 12390
rect 9646 12362 9674 12367
rect 9254 11923 9282 11942
rect 9366 12361 9674 12362
rect 9366 12335 9647 12361
rect 9673 12335 9674 12361
rect 9366 12334 9674 12335
rect 9366 11969 9394 12334
rect 9646 12329 9674 12334
rect 9702 12138 9730 12446
rect 9758 12473 9786 12614
rect 9758 12447 9759 12473
rect 9785 12447 9786 12473
rect 9758 12441 9786 12447
rect 9814 12418 9842 12782
rect 10038 12753 10066 12782
rect 10038 12727 10039 12753
rect 10065 12727 10066 12753
rect 10038 12721 10066 12727
rect 10094 12753 10122 12759
rect 10094 12727 10095 12753
rect 10121 12727 10122 12753
rect 9870 12698 9898 12703
rect 9982 12698 10010 12703
rect 9898 12670 9954 12698
rect 9870 12665 9898 12670
rect 9926 12641 9954 12670
rect 9982 12651 10010 12670
rect 9926 12615 9927 12641
rect 9953 12615 9954 12641
rect 9926 12609 9954 12615
rect 10094 12642 10122 12727
rect 10094 12609 10122 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12385 9842 12390
rect 9982 12361 10010 12367
rect 9982 12335 9983 12361
rect 10009 12335 10010 12361
rect 9814 12250 9842 12255
rect 9814 12203 9842 12222
rect 9982 12138 10010 12335
rect 10150 12362 10178 12782
rect 10206 12754 10234 13063
rect 10262 13593 10402 13594
rect 10262 13567 10375 13593
rect 10401 13567 10402 13593
rect 10262 13566 10402 13567
rect 10262 12865 10290 13566
rect 10374 13561 10402 13566
rect 11774 13537 11802 13543
rect 11774 13511 11775 13537
rect 11801 13511 11802 13537
rect 10710 13426 10738 13431
rect 10654 13425 10738 13426
rect 10654 13399 10711 13425
rect 10737 13399 10738 13425
rect 10654 13398 10738 13399
rect 10318 13202 10346 13207
rect 10430 13202 10458 13207
rect 10654 13202 10682 13398
rect 10710 13393 10738 13398
rect 10878 13202 10906 13207
rect 10346 13201 10682 13202
rect 10346 13175 10431 13201
rect 10457 13175 10682 13201
rect 10346 13174 10682 13175
rect 10822 13174 10878 13202
rect 10318 13169 10346 13174
rect 10430 13169 10458 13174
rect 10710 13146 10738 13151
rect 10710 13099 10738 13118
rect 10262 12839 10263 12865
rect 10289 12839 10290 12865
rect 10262 12833 10290 12839
rect 10710 12866 10738 12871
rect 10710 12809 10738 12838
rect 10710 12783 10711 12809
rect 10737 12783 10738 12809
rect 10710 12777 10738 12783
rect 10822 12810 10850 13174
rect 10878 13169 10906 13174
rect 11774 13146 11802 13511
rect 11774 13113 11802 13118
rect 11046 13090 11074 13095
rect 12054 13090 12082 15946
rect 13174 13594 13202 18606
rect 13006 13593 13202 13594
rect 13006 13567 13175 13593
rect 13201 13567 13202 13593
rect 13006 13566 13202 13567
rect 12110 13481 12138 13487
rect 12110 13455 12111 13481
rect 12137 13455 12138 13481
rect 12110 13258 12138 13455
rect 12110 13225 12138 13230
rect 12334 13482 12362 13487
rect 13006 13454 13034 13566
rect 13174 13561 13202 13566
rect 12334 13146 12362 13454
rect 12950 13426 13034 13454
rect 13398 13482 13426 13487
rect 13426 13454 13482 13482
rect 13398 13435 13426 13454
rect 12670 13258 12698 13263
rect 12670 13211 12698 13230
rect 12726 13202 12754 13207
rect 12726 13155 12754 13174
rect 12950 13146 12978 13426
rect 13118 13258 13146 13263
rect 13118 13211 13146 13230
rect 12334 13099 12362 13118
rect 12894 13145 12978 13146
rect 12894 13119 12951 13145
rect 12977 13119 12978 13145
rect 12894 13118 12978 13119
rect 12110 13090 12138 13095
rect 11046 13089 11298 13090
rect 11046 13063 11047 13089
rect 11073 13063 11298 13089
rect 11046 13062 11298 13063
rect 12054 13089 12138 13090
rect 12054 13063 12111 13089
rect 12137 13063 12138 13089
rect 12054 13062 12138 13063
rect 11046 13057 11074 13062
rect 10206 12721 10234 12726
rect 10654 12698 10682 12703
rect 10654 12651 10682 12670
rect 10766 12642 10794 12647
rect 10766 12595 10794 12614
rect 10206 12474 10234 12479
rect 10234 12446 10290 12474
rect 10206 12441 10234 12446
rect 10262 12417 10290 12446
rect 10262 12391 10263 12417
rect 10289 12391 10290 12417
rect 10262 12385 10290 12391
rect 10206 12362 10234 12367
rect 10150 12361 10234 12362
rect 10150 12335 10207 12361
rect 10233 12335 10234 12361
rect 10150 12334 10234 12335
rect 10206 12329 10234 12334
rect 10318 12334 10626 12362
rect 10094 12250 10122 12255
rect 10318 12250 10346 12334
rect 10094 12249 10346 12250
rect 10094 12223 10095 12249
rect 10121 12223 10346 12249
rect 10094 12222 10346 12223
rect 10486 12250 10514 12255
rect 10094 12217 10122 12222
rect 9702 12110 10010 12138
rect 10430 12082 10458 12087
rect 9366 11943 9367 11969
rect 9393 11943 9394 11969
rect 9366 11690 9394 11943
rect 9534 12025 9562 12031
rect 9534 11999 9535 12025
rect 9561 11999 9562 12025
rect 9534 11914 9562 11999
rect 9534 11881 9562 11886
rect 9814 11913 9842 11919
rect 9814 11887 9815 11913
rect 9841 11887 9842 11913
rect 9590 11858 9618 11863
rect 9366 11689 9506 11690
rect 9366 11663 9367 11689
rect 9393 11663 9506 11689
rect 9366 11662 9506 11663
rect 9366 11657 9394 11662
rect 9198 11215 9199 11241
rect 9225 11215 9226 11241
rect 9198 10122 9226 11215
rect 9478 11129 9506 11662
rect 9534 11634 9562 11639
rect 9534 11587 9562 11606
rect 9534 11242 9562 11247
rect 9534 11185 9562 11214
rect 9534 11159 9535 11185
rect 9561 11159 9562 11185
rect 9534 11153 9562 11159
rect 9478 11103 9479 11129
rect 9505 11103 9506 11129
rect 9310 10906 9338 10911
rect 9254 10850 9282 10855
rect 9254 10803 9282 10822
rect 9254 10570 9282 10575
rect 9254 10401 9282 10542
rect 9254 10375 9255 10401
rect 9281 10375 9282 10401
rect 9254 10369 9282 10375
rect 9310 10290 9338 10878
rect 9478 10457 9506 11103
rect 9478 10431 9479 10457
rect 9505 10431 9506 10457
rect 9478 10425 9506 10431
rect 9534 11074 9562 11079
rect 9590 11074 9618 11830
rect 9814 11858 9842 11887
rect 9870 11914 9898 11919
rect 9870 11867 9898 11886
rect 9814 11825 9842 11830
rect 9982 11858 10010 11877
rect 9982 11825 10010 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11746 10122 11751
rect 9814 11633 9842 11639
rect 9814 11607 9815 11633
rect 9841 11607 9842 11633
rect 9758 11522 9786 11527
rect 9702 11466 9730 11471
rect 9562 11046 9618 11074
rect 9646 11465 9730 11466
rect 9646 11439 9703 11465
rect 9729 11439 9730 11465
rect 9646 11438 9730 11439
rect 9030 10121 9114 10122
rect 9030 10095 9031 10121
rect 9057 10095 9114 10121
rect 9030 10094 9114 10095
rect 9030 10089 9058 10094
rect 8806 10065 8834 10071
rect 8806 10039 8807 10065
rect 8833 10039 8834 10065
rect 8806 9898 8834 10039
rect 8806 9865 8834 9870
rect 8918 10010 8946 10015
rect 8862 9730 8890 9735
rect 8862 9618 8890 9702
rect 8862 9585 8890 9590
rect 8806 9562 8834 9567
rect 8806 9515 8834 9534
rect 8862 9506 8890 9511
rect 8918 9506 8946 9982
rect 8974 9954 9002 9959
rect 8974 9907 9002 9926
rect 9086 9673 9114 10094
rect 9198 10089 9226 10094
rect 9254 10262 9338 10290
rect 9254 9954 9282 10262
rect 9366 10065 9394 10071
rect 9366 10039 9367 10065
rect 9393 10039 9394 10065
rect 9366 10010 9394 10039
rect 9366 9977 9394 9982
rect 9478 10009 9506 10015
rect 9478 9983 9479 10009
rect 9505 9983 9506 10009
rect 9198 9926 9282 9954
rect 9310 9954 9338 9959
rect 9198 9786 9226 9926
rect 9198 9758 9282 9786
rect 9086 9647 9087 9673
rect 9113 9647 9114 9673
rect 9086 9641 9114 9647
rect 9254 9673 9282 9758
rect 9254 9647 9255 9673
rect 9281 9647 9282 9673
rect 9254 9641 9282 9647
rect 8862 9505 8946 9506
rect 8862 9479 8863 9505
rect 8889 9479 8946 9505
rect 8862 9478 8946 9479
rect 9142 9618 9170 9623
rect 8862 9282 8890 9478
rect 8862 9249 8890 9254
rect 9030 9450 9058 9455
rect 8806 8834 8834 8839
rect 8750 8806 8806 8834
rect 8806 8787 8834 8806
rect 8974 8442 9002 8447
rect 8750 8106 8778 8111
rect 8974 8106 9002 8414
rect 8750 8105 9002 8106
rect 8750 8079 8751 8105
rect 8777 8079 9002 8105
rect 8750 8078 9002 8079
rect 8750 8073 8778 8078
rect 8302 8023 8303 8049
rect 8329 8023 8330 8049
rect 8302 8017 8330 8023
rect 8526 8049 8554 8055
rect 8526 8023 8527 8049
rect 8553 8023 8554 8049
rect 6902 7686 7322 7714
rect 8302 7938 8330 7943
rect 6902 7657 6930 7686
rect 6902 7631 6903 7657
rect 6929 7631 6930 7657
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 6846 7266 6874 7271
rect 6902 7266 6930 7631
rect 8302 7658 8330 7910
rect 8358 7937 8386 7943
rect 8358 7911 8359 7937
rect 8385 7911 8386 7937
rect 8358 7826 8386 7911
rect 8414 7938 8442 7943
rect 8526 7938 8554 8023
rect 8974 8049 9002 8078
rect 8974 8023 8975 8049
rect 9001 8023 9002 8049
rect 8974 8017 9002 8023
rect 9030 8049 9058 9422
rect 9030 8023 9031 8049
rect 9057 8023 9058 8049
rect 8694 7938 8722 7943
rect 9030 7938 9058 8023
rect 9086 8050 9114 8055
rect 9142 8050 9170 9590
rect 9310 9281 9338 9926
rect 9422 9954 9450 9959
rect 9422 9907 9450 9926
rect 9310 9255 9311 9281
rect 9337 9255 9338 9281
rect 9310 9249 9338 9255
rect 9366 9282 9394 9287
rect 9366 9281 9450 9282
rect 9366 9255 9367 9281
rect 9393 9255 9450 9281
rect 9366 9254 9450 9255
rect 9366 9249 9394 9254
rect 9366 9114 9394 9119
rect 9198 9113 9394 9114
rect 9198 9087 9367 9113
rect 9393 9087 9394 9113
rect 9198 9086 9394 9087
rect 9198 8889 9226 9086
rect 9366 9081 9394 9086
rect 9422 9114 9450 9254
rect 9422 9081 9450 9086
rect 9198 8863 9199 8889
rect 9225 8863 9226 8889
rect 9198 8857 9226 8863
rect 9478 8778 9506 9983
rect 9534 9170 9562 11046
rect 9646 10906 9674 11438
rect 9702 11433 9730 11438
rect 9702 11186 9730 11191
rect 9702 11139 9730 11158
rect 9646 10873 9674 10878
rect 9758 10401 9786 11494
rect 9814 10570 9842 11607
rect 9982 11129 10010 11135
rect 9982 11103 9983 11129
rect 10009 11103 10010 11129
rect 9982 11074 10010 11103
rect 9982 11041 10010 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10094 10906 10122 11718
rect 10430 11689 10458 12054
rect 10430 11663 10431 11689
rect 10457 11663 10458 11689
rect 10430 11657 10458 11663
rect 10318 11633 10346 11639
rect 10318 11607 10319 11633
rect 10345 11607 10346 11633
rect 10262 11577 10290 11583
rect 10262 11551 10263 11577
rect 10289 11551 10290 11577
rect 10262 11522 10290 11551
rect 10262 11489 10290 11494
rect 9814 10537 9842 10542
rect 10038 10878 10122 10906
rect 10038 10513 10066 10878
rect 10318 10626 10346 11607
rect 10262 10598 10346 10626
rect 10374 11186 10402 11191
rect 10038 10487 10039 10513
rect 10065 10487 10066 10513
rect 10038 10481 10066 10487
rect 10150 10570 10178 10575
rect 9758 10375 9759 10401
rect 9785 10375 9786 10401
rect 9758 10369 9786 10375
rect 9814 10374 10010 10402
rect 9758 10066 9786 10071
rect 9814 10066 9842 10374
rect 9982 10345 10010 10374
rect 9982 10319 9983 10345
rect 10009 10319 10010 10345
rect 9982 10313 10010 10319
rect 10150 10345 10178 10542
rect 10262 10402 10290 10598
rect 10318 10514 10346 10519
rect 10374 10514 10402 11158
rect 10486 11018 10514 12222
rect 10542 11633 10570 11639
rect 10542 11607 10543 11633
rect 10569 11607 10570 11633
rect 10542 11578 10570 11607
rect 10542 11186 10570 11550
rect 10598 11522 10626 12334
rect 10766 12026 10794 12031
rect 10822 12026 10850 12782
rect 11270 12809 11298 13062
rect 11550 12866 11578 12871
rect 11270 12783 11271 12809
rect 11297 12783 11298 12809
rect 11270 12777 11298 12783
rect 11382 12865 11578 12866
rect 11382 12839 11551 12865
rect 11577 12839 11578 12865
rect 11382 12838 11578 12839
rect 11102 12753 11130 12759
rect 11102 12727 11103 12753
rect 11129 12727 11130 12753
rect 11102 12642 11130 12727
rect 11382 12753 11410 12838
rect 11550 12833 11578 12838
rect 11382 12727 11383 12753
rect 11409 12727 11410 12753
rect 11382 12721 11410 12727
rect 11830 12754 11858 12759
rect 11102 12081 11130 12614
rect 11102 12055 11103 12081
rect 11129 12055 11130 12081
rect 11102 12049 11130 12055
rect 11158 12697 11186 12703
rect 11158 12671 11159 12697
rect 11185 12671 11186 12697
rect 10766 12025 10850 12026
rect 10766 11999 10767 12025
rect 10793 11999 10850 12025
rect 10766 11998 10850 11999
rect 10766 11993 10794 11998
rect 11046 11970 11074 11975
rect 11158 11970 11186 12671
rect 11494 12697 11522 12703
rect 11494 12671 11495 12697
rect 11521 12671 11522 12697
rect 11494 12082 11522 12671
rect 11550 12698 11578 12703
rect 11550 12651 11578 12670
rect 11774 12642 11802 12647
rect 11494 12049 11522 12054
rect 11718 12614 11774 12642
rect 11438 11970 11466 11975
rect 11718 11970 11746 12614
rect 11774 12609 11802 12614
rect 11046 11969 11130 11970
rect 11046 11943 11047 11969
rect 11073 11943 11130 11969
rect 11046 11942 11130 11943
rect 11046 11937 11074 11942
rect 10766 11914 10794 11919
rect 10710 11857 10738 11863
rect 10710 11831 10711 11857
rect 10737 11831 10738 11857
rect 10654 11746 10682 11751
rect 10654 11689 10682 11718
rect 10654 11663 10655 11689
rect 10681 11663 10682 11689
rect 10654 11657 10682 11663
rect 10654 11522 10682 11527
rect 10598 11521 10682 11522
rect 10598 11495 10655 11521
rect 10681 11495 10682 11521
rect 10598 11494 10682 11495
rect 10542 11153 10570 11158
rect 10598 11298 10626 11303
rect 10598 11074 10626 11270
rect 10654 11186 10682 11494
rect 10710 11522 10738 11831
rect 10710 11489 10738 11494
rect 10766 11577 10794 11886
rect 10822 11858 10850 11863
rect 10822 11811 10850 11830
rect 10766 11551 10767 11577
rect 10793 11551 10794 11577
rect 10654 11158 10738 11186
rect 10654 11074 10682 11079
rect 10598 11073 10682 11074
rect 10598 11047 10655 11073
rect 10681 11047 10682 11073
rect 10598 11046 10682 11047
rect 10654 11041 10682 11046
rect 10486 10990 10626 11018
rect 10598 10962 10626 10990
rect 10598 10934 10682 10962
rect 10318 10513 10402 10514
rect 10318 10487 10319 10513
rect 10345 10487 10402 10513
rect 10318 10486 10402 10487
rect 10598 10850 10626 10855
rect 10318 10481 10346 10486
rect 10374 10402 10402 10407
rect 10262 10401 10402 10402
rect 10262 10375 10375 10401
rect 10401 10375 10402 10401
rect 10262 10374 10402 10375
rect 10150 10319 10151 10345
rect 10177 10319 10178 10345
rect 10150 10313 10178 10319
rect 9870 10290 9898 10309
rect 9870 10257 9898 10262
rect 10262 10289 10290 10295
rect 10262 10263 10263 10289
rect 10289 10263 10290 10289
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9786 10038 9842 10066
rect 9702 10010 9730 10015
rect 9590 10009 9730 10010
rect 9590 9983 9703 10009
rect 9729 9983 9730 10009
rect 9590 9982 9730 9983
rect 9590 9673 9618 9982
rect 9702 9977 9730 9982
rect 9590 9647 9591 9673
rect 9617 9647 9618 9673
rect 9590 9506 9618 9647
rect 9758 9618 9786 10038
rect 10262 9730 10290 10263
rect 10094 9702 10290 9730
rect 10374 10010 10402 10374
rect 9982 9674 10010 9679
rect 9758 9585 9786 9590
rect 9814 9673 10010 9674
rect 9814 9647 9983 9673
rect 10009 9647 10010 9673
rect 9814 9646 10010 9647
rect 9590 9473 9618 9478
rect 9702 9561 9730 9567
rect 9702 9535 9703 9561
rect 9729 9535 9730 9561
rect 9590 9170 9618 9175
rect 9534 9142 9590 9170
rect 9590 9123 9618 9142
rect 9702 9170 9730 9535
rect 9758 9505 9786 9511
rect 9758 9479 9759 9505
rect 9785 9479 9786 9505
rect 9758 9226 9786 9479
rect 9758 9193 9786 9198
rect 9702 9137 9730 9142
rect 9478 8745 9506 8750
rect 9814 8442 9842 9646
rect 9982 9641 10010 9646
rect 10038 9618 10066 9623
rect 10094 9618 10122 9702
rect 10038 9617 10122 9618
rect 10038 9591 10039 9617
rect 10065 9591 10122 9617
rect 10038 9590 10122 9591
rect 10206 9618 10234 9623
rect 9926 9562 9954 9567
rect 9926 9515 9954 9534
rect 10038 9506 10066 9590
rect 10206 9571 10234 9590
rect 10038 9473 10066 9478
rect 10150 9562 10178 9567
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9870 9226 9898 9231
rect 9870 9179 9898 9198
rect 10150 9225 10178 9534
rect 10150 9199 10151 9225
rect 10177 9199 10178 9225
rect 10150 9193 10178 9199
rect 10206 9170 10234 9175
rect 10206 8890 10234 9142
rect 10374 9113 10402 9982
rect 10598 9954 10626 10822
rect 10654 10513 10682 10934
rect 10654 10487 10655 10513
rect 10681 10487 10682 10513
rect 10654 10481 10682 10487
rect 10710 10458 10738 11158
rect 10766 11185 10794 11551
rect 10990 11578 11018 11583
rect 11102 11578 11130 11942
rect 11158 11937 11186 11942
rect 11214 11969 11746 11970
rect 11214 11943 11439 11969
rect 11465 11943 11746 11969
rect 11214 11942 11746 11943
rect 11158 11858 11186 11863
rect 11158 11811 11186 11830
rect 11158 11690 11186 11695
rect 11214 11690 11242 11942
rect 11438 11937 11466 11942
rect 11158 11689 11242 11690
rect 11158 11663 11159 11689
rect 11185 11663 11242 11689
rect 11158 11662 11242 11663
rect 11270 11857 11298 11863
rect 11270 11831 11271 11857
rect 11297 11831 11298 11857
rect 11158 11657 11186 11662
rect 11270 11578 11298 11831
rect 11018 11550 11074 11578
rect 11102 11550 11298 11578
rect 10990 11531 11018 11550
rect 10766 11159 10767 11185
rect 10793 11159 10794 11185
rect 10766 10850 10794 11159
rect 11046 11185 11074 11550
rect 11046 11159 11047 11185
rect 11073 11159 11074 11185
rect 11046 11153 11074 11159
rect 11102 11185 11130 11191
rect 11102 11159 11103 11185
rect 11129 11159 11130 11185
rect 10822 11130 10850 11135
rect 10990 11130 11018 11135
rect 10850 11102 10906 11130
rect 10822 11097 10850 11102
rect 10766 10817 10794 10822
rect 10878 10458 10906 11102
rect 10990 11083 11018 11102
rect 11102 10514 11130 11159
rect 11270 10906 11298 11550
rect 11326 11746 11354 11751
rect 11326 11185 11354 11718
rect 11718 11690 11746 11942
rect 11774 11690 11802 11695
rect 11718 11689 11802 11690
rect 11718 11663 11775 11689
rect 11801 11663 11802 11689
rect 11718 11662 11802 11663
rect 11774 11657 11802 11662
rect 11326 11159 11327 11185
rect 11353 11159 11354 11185
rect 11326 11153 11354 11159
rect 11494 11634 11522 11639
rect 11494 11130 11522 11606
rect 11830 11634 11858 12726
rect 12110 12698 12138 13062
rect 12614 13033 12642 13039
rect 12614 13007 12615 13033
rect 12641 13007 12642 13033
rect 12614 12865 12642 13007
rect 12614 12839 12615 12865
rect 12641 12839 12642 12865
rect 12614 12833 12642 12839
rect 12334 12754 12362 12759
rect 12334 12707 12362 12726
rect 12110 12665 12138 12670
rect 12278 12697 12306 12703
rect 12278 12671 12279 12697
rect 12305 12671 12306 12697
rect 12278 12642 12306 12671
rect 12390 12698 12418 12703
rect 12390 12651 12418 12670
rect 12782 12697 12810 12703
rect 12782 12671 12783 12697
rect 12809 12671 12810 12697
rect 12278 12609 12306 12614
rect 12782 12306 12810 12671
rect 12838 12698 12866 12703
rect 12894 12698 12922 13118
rect 12950 13113 12978 13118
rect 13454 13146 13482 13454
rect 14294 13258 14322 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 14294 13225 14322 13230
rect 18942 13537 18970 13543
rect 18942 13511 18943 13537
rect 18969 13511 18970 13537
rect 13454 13145 13706 13146
rect 13454 13119 13455 13145
rect 13481 13119 13706 13145
rect 13454 13118 13706 13119
rect 13454 13113 13482 13118
rect 12838 12697 12922 12698
rect 12838 12671 12839 12697
rect 12865 12671 12922 12697
rect 12838 12670 12922 12671
rect 12950 12698 12978 12703
rect 12838 12665 12866 12670
rect 12950 12651 12978 12670
rect 13678 12474 13706 13118
rect 18830 13145 18858 13151
rect 18830 13119 18831 13145
rect 18857 13119 18858 13145
rect 13790 13089 13818 13095
rect 13790 13063 13791 13089
rect 13817 13063 13818 13089
rect 13734 12866 13762 12871
rect 13790 12866 13818 13063
rect 13734 12865 13818 12866
rect 13734 12839 13735 12865
rect 13761 12839 13818 12865
rect 13734 12838 13818 12839
rect 14854 13089 14882 13095
rect 14854 13063 14855 13089
rect 14881 13063 14882 13089
rect 13734 12833 13762 12838
rect 14294 12782 14770 12810
rect 14238 12754 14266 12759
rect 13790 12698 13818 12703
rect 13790 12651 13818 12670
rect 14238 12697 14266 12726
rect 14294 12753 14322 12782
rect 14294 12727 14295 12753
rect 14321 12727 14322 12753
rect 14294 12721 14322 12727
rect 14742 12754 14770 12782
rect 14798 12754 14826 12759
rect 14742 12753 14826 12754
rect 14742 12727 14799 12753
rect 14825 12727 14826 12753
rect 14742 12726 14826 12727
rect 14798 12721 14826 12726
rect 14238 12671 14239 12697
rect 14265 12671 14266 12697
rect 14238 12665 14266 12671
rect 14518 12698 14546 12703
rect 14518 12651 14546 12670
rect 14630 12698 14658 12703
rect 14630 12651 14658 12670
rect 14686 12697 14714 12703
rect 14686 12671 14687 12697
rect 14713 12671 14714 12697
rect 13734 12642 13762 12647
rect 13734 12595 13762 12614
rect 14126 12642 14154 12647
rect 14126 12641 14210 12642
rect 14126 12615 14127 12641
rect 14153 12615 14210 12641
rect 14126 12614 14210 12615
rect 14126 12609 14154 12614
rect 13678 12473 13874 12474
rect 13678 12447 13679 12473
rect 13705 12447 13874 12473
rect 13678 12446 13874 12447
rect 13678 12441 13706 12446
rect 12782 11689 12810 12278
rect 13846 12361 13874 12446
rect 14182 12418 14210 12614
rect 14686 12586 14714 12671
rect 14854 12698 14882 13063
rect 15078 13089 15106 13095
rect 15078 13063 15079 13089
rect 15105 13063 15106 13089
rect 14854 12665 14882 12670
rect 14910 13034 14938 13039
rect 14910 12697 14938 13006
rect 14910 12671 14911 12697
rect 14937 12671 14938 12697
rect 14910 12665 14938 12671
rect 14966 12697 14994 12703
rect 14966 12671 14967 12697
rect 14993 12671 14994 12697
rect 14966 12586 14994 12671
rect 14686 12558 14994 12586
rect 14238 12418 14266 12423
rect 14182 12417 14266 12418
rect 14182 12391 14239 12417
rect 14265 12391 14266 12417
rect 14182 12390 14266 12391
rect 14238 12385 14266 12390
rect 13846 12335 13847 12361
rect 13873 12335 13874 12361
rect 13846 12026 13874 12335
rect 13846 11993 13874 11998
rect 14014 12026 14042 12031
rect 12782 11663 12783 11689
rect 12809 11663 12810 11689
rect 12782 11657 12810 11663
rect 11830 11587 11858 11606
rect 13342 11633 13370 11639
rect 13342 11607 13343 11633
rect 13369 11607 13370 11633
rect 11662 11578 11690 11583
rect 12054 11578 12082 11583
rect 11662 11577 11746 11578
rect 11662 11551 11663 11577
rect 11689 11551 11746 11577
rect 11662 11550 11746 11551
rect 11662 11545 11690 11550
rect 11494 11083 11522 11102
rect 11298 10878 11410 10906
rect 11270 10873 11298 10878
rect 11326 10793 11354 10799
rect 11326 10767 11327 10793
rect 11353 10767 11354 10793
rect 11046 10486 11130 10514
rect 11214 10514 11242 10519
rect 10934 10458 10962 10463
rect 10710 10430 10794 10458
rect 10598 9338 10626 9926
rect 10710 10346 10738 10351
rect 10710 9561 10738 10318
rect 10710 9535 10711 9561
rect 10737 9535 10738 9561
rect 10710 9529 10738 9535
rect 10598 9305 10626 9310
rect 10654 9225 10682 9231
rect 10654 9199 10655 9225
rect 10681 9199 10682 9225
rect 10654 9170 10682 9199
rect 10654 9137 10682 9142
rect 10374 9087 10375 9113
rect 10401 9087 10402 9113
rect 10374 9081 10402 9087
rect 10262 8890 10290 8895
rect 10206 8889 10290 8890
rect 10206 8863 10263 8889
rect 10289 8863 10290 8889
rect 10206 8862 10290 8863
rect 10262 8857 10290 8862
rect 10710 8834 10738 8839
rect 10710 8787 10738 8806
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9814 8395 9842 8414
rect 9926 8498 9954 8503
rect 9086 8049 9170 8050
rect 9086 8023 9087 8049
rect 9113 8023 9170 8049
rect 9086 8022 9170 8023
rect 9086 8017 9114 8022
rect 8526 7910 8694 7938
rect 8414 7891 8442 7910
rect 8694 7891 8722 7910
rect 8750 7910 9058 7938
rect 9254 7938 9282 7943
rect 8358 7798 8442 7826
rect 7182 7602 7210 7607
rect 7182 7321 7210 7574
rect 7238 7601 7266 7607
rect 7238 7575 7239 7601
rect 7265 7575 7266 7601
rect 7238 7378 7266 7575
rect 8302 7601 8330 7630
rect 8302 7575 8303 7601
rect 8329 7575 8330 7601
rect 8302 7569 8330 7575
rect 7238 7345 7266 7350
rect 8414 7377 8442 7798
rect 8694 7714 8722 7719
rect 8750 7714 8778 7910
rect 9086 7770 9114 7775
rect 8694 7713 8778 7714
rect 8694 7687 8695 7713
rect 8721 7687 8778 7713
rect 8694 7686 8778 7687
rect 8862 7769 9114 7770
rect 8862 7743 9087 7769
rect 9113 7743 9114 7769
rect 8862 7742 9114 7743
rect 8862 7713 8890 7742
rect 9086 7737 9114 7742
rect 8862 7687 8863 7713
rect 8889 7687 8890 7713
rect 8694 7681 8722 7686
rect 8862 7681 8890 7687
rect 9198 7713 9226 7719
rect 9198 7687 9199 7713
rect 9225 7687 9226 7713
rect 8638 7658 8666 7663
rect 8414 7351 8415 7377
rect 8441 7351 8442 7377
rect 8414 7345 8442 7351
rect 8470 7378 8498 7383
rect 7182 7295 7183 7321
rect 7209 7295 7210 7321
rect 7182 7289 7210 7295
rect 8246 7322 8274 7327
rect 8246 7275 8274 7294
rect 8470 7321 8498 7350
rect 8470 7295 8471 7321
rect 8497 7295 8498 7321
rect 8470 7289 8498 7295
rect 8582 7378 8610 7383
rect 6846 7265 6902 7266
rect 6846 7239 6847 7265
rect 6873 7239 6902 7265
rect 6846 7238 6902 7239
rect 6846 7233 6874 7238
rect 6902 7219 6930 7238
rect 8358 7266 8386 7271
rect 8358 6986 8386 7238
rect 8582 7265 8610 7350
rect 8582 7239 8583 7265
rect 8609 7239 8610 7265
rect 8582 7233 8610 7239
rect 8358 6985 8610 6986
rect 8358 6959 8359 6985
rect 8385 6959 8610 6985
rect 8358 6958 8610 6959
rect 8358 6953 8386 6958
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 8582 6481 8610 6958
rect 8582 6455 8583 6481
rect 8609 6455 8610 6481
rect 8582 6449 8610 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8078 2114 8106 2119
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8078 400 8106 2086
rect 8638 1777 8666 7630
rect 8974 7657 9002 7663
rect 8974 7631 8975 7657
rect 9001 7631 9002 7657
rect 8750 7602 8778 7621
rect 8750 7569 8778 7574
rect 8974 7378 9002 7631
rect 9198 7378 9226 7687
rect 9254 7713 9282 7910
rect 9254 7687 9255 7713
rect 9281 7687 9282 7713
rect 9254 7681 9282 7687
rect 9310 7937 9338 7943
rect 9926 7938 9954 8470
rect 9310 7911 9311 7937
rect 9337 7911 9338 7937
rect 9310 7574 9338 7911
rect 9814 7910 9954 7938
rect 9814 7574 9842 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9310 7546 9450 7574
rect 9814 7546 9954 7574
rect 8974 7345 9002 7350
rect 9086 7350 9226 7378
rect 9310 7378 9338 7383
rect 8694 7322 8722 7327
rect 8694 2169 8722 7294
rect 9086 7322 9114 7350
rect 9310 7331 9338 7350
rect 9422 7377 9450 7546
rect 9422 7351 9423 7377
rect 9449 7351 9450 7377
rect 9422 7345 9450 7351
rect 9926 7378 9954 7546
rect 9926 7377 10234 7378
rect 9926 7351 9927 7377
rect 9953 7351 10234 7377
rect 9926 7350 10234 7351
rect 9926 7345 9954 7350
rect 9086 7289 9114 7294
rect 9758 7321 9786 7327
rect 9758 7295 9759 7321
rect 9785 7295 9786 7321
rect 8806 7266 8834 7271
rect 8806 7219 8834 7238
rect 9310 7266 9338 7271
rect 8974 7210 9002 7215
rect 8974 6537 9002 7182
rect 9254 7210 9282 7215
rect 9254 7163 9282 7182
rect 9310 6874 9338 7238
rect 9534 7266 9562 7271
rect 9758 7266 9786 7295
rect 9534 7265 9786 7266
rect 9534 7239 9535 7265
rect 9561 7239 9786 7265
rect 9534 7238 9786 7239
rect 10206 7266 10234 7350
rect 10766 7377 10794 10430
rect 10878 10457 10962 10458
rect 10878 10431 10935 10457
rect 10961 10431 10962 10457
rect 10878 10430 10962 10431
rect 10822 10401 10850 10407
rect 10822 10375 10823 10401
rect 10849 10375 10850 10401
rect 10822 10066 10850 10375
rect 10878 10346 10906 10430
rect 10934 10425 10962 10430
rect 10878 10313 10906 10318
rect 10850 10038 10906 10066
rect 10822 10033 10850 10038
rect 10878 9618 10906 10038
rect 10822 9338 10850 9343
rect 10878 9338 10906 9590
rect 10934 9561 10962 9567
rect 10934 9535 10935 9561
rect 10961 9535 10962 9561
rect 10934 9506 10962 9535
rect 10934 9473 10962 9478
rect 10822 9337 10906 9338
rect 10822 9311 10823 9337
rect 10849 9311 10906 9337
rect 10822 9310 10906 9311
rect 10822 9305 10850 9310
rect 10990 9226 11018 9231
rect 10990 9179 11018 9198
rect 11046 8498 11074 10486
rect 11102 10401 11130 10407
rect 11102 10375 11103 10401
rect 11129 10375 11130 10401
rect 11102 10290 11130 10375
rect 11214 10401 11242 10486
rect 11214 10375 11215 10401
rect 11241 10375 11242 10401
rect 11214 10369 11242 10375
rect 11326 10402 11354 10767
rect 11326 10369 11354 10374
rect 11102 9618 11130 10262
rect 11158 10289 11186 10295
rect 11158 10263 11159 10289
rect 11185 10263 11186 10289
rect 11158 10010 11186 10263
rect 11158 9977 11186 9982
rect 11158 9618 11186 9623
rect 11102 9617 11242 9618
rect 11102 9591 11159 9617
rect 11185 9591 11242 9617
rect 11102 9590 11242 9591
rect 11158 9585 11186 9590
rect 11214 9562 11242 9590
rect 11214 9169 11242 9534
rect 11270 9562 11298 9567
rect 11270 9561 11354 9562
rect 11270 9535 11271 9561
rect 11297 9535 11354 9561
rect 11270 9534 11354 9535
rect 11270 9529 11298 9534
rect 11214 9143 11215 9169
rect 11241 9143 11242 9169
rect 11214 9137 11242 9143
rect 11326 8890 11354 9534
rect 11326 8777 11354 8862
rect 11382 8834 11410 10878
rect 11550 10849 11578 10855
rect 11550 10823 11551 10849
rect 11577 10823 11578 10849
rect 11494 10793 11522 10799
rect 11494 10767 11495 10793
rect 11521 10767 11522 10793
rect 11494 10066 11522 10767
rect 11550 10514 11578 10823
rect 11662 10794 11690 10799
rect 11662 10747 11690 10766
rect 11550 10481 11578 10486
rect 11438 10038 11494 10066
rect 11438 9617 11466 10038
rect 11494 10033 11522 10038
rect 11662 10402 11690 10407
rect 11662 10065 11690 10374
rect 11662 10039 11663 10065
rect 11689 10039 11690 10065
rect 11662 10033 11690 10039
rect 11438 9591 11439 9617
rect 11465 9591 11466 9617
rect 11438 9585 11466 9591
rect 11550 9898 11578 9903
rect 11550 9505 11578 9870
rect 11550 9479 11551 9505
rect 11577 9479 11578 9505
rect 11550 9450 11578 9479
rect 11550 9417 11578 9422
rect 11662 9506 11690 9511
rect 11494 9281 11522 9287
rect 11494 9255 11495 9281
rect 11521 9255 11522 9281
rect 11494 9114 11522 9255
rect 11494 8834 11522 9086
rect 11662 9225 11690 9478
rect 11662 9199 11663 9225
rect 11689 9199 11690 9225
rect 11382 8833 11466 8834
rect 11382 8807 11383 8833
rect 11409 8807 11466 8833
rect 11382 8806 11466 8807
rect 11382 8801 11410 8806
rect 11326 8751 11327 8777
rect 11353 8751 11354 8777
rect 11326 8745 11354 8751
rect 11214 8722 11242 8727
rect 11438 8722 11466 8806
rect 11494 8801 11522 8806
rect 11606 8834 11634 8839
rect 11662 8834 11690 9199
rect 11606 8833 11690 8834
rect 11606 8807 11607 8833
rect 11633 8807 11690 8833
rect 11606 8806 11690 8807
rect 11606 8801 11634 8806
rect 11662 8722 11690 8727
rect 11214 8721 11298 8722
rect 11214 8695 11215 8721
rect 11241 8695 11298 8721
rect 11214 8694 11298 8695
rect 11438 8721 11690 8722
rect 11438 8695 11663 8721
rect 11689 8695 11690 8721
rect 11438 8694 11690 8695
rect 11214 8689 11242 8694
rect 11046 8465 11074 8470
rect 10822 7713 10850 7719
rect 10822 7687 10823 7713
rect 10849 7687 10850 7713
rect 10822 7574 10850 7687
rect 10990 7714 11018 7719
rect 11270 7714 11298 8694
rect 11662 8689 11690 8694
rect 11718 8050 11746 11550
rect 11998 11242 12026 11247
rect 11998 11185 12026 11214
rect 11998 11159 11999 11185
rect 12025 11159 12026 11185
rect 11998 11153 12026 11159
rect 12054 11129 12082 11550
rect 12670 11577 12698 11583
rect 12670 11551 12671 11577
rect 12697 11551 12698 11577
rect 12054 11103 12055 11129
rect 12081 11103 12082 11129
rect 11942 10906 11970 10911
rect 11942 10859 11970 10878
rect 12054 10458 12082 11103
rect 12390 11185 12418 11191
rect 12390 11159 12391 11185
rect 12417 11159 12418 11185
rect 12166 11074 12194 11079
rect 12166 11027 12194 11046
rect 12390 10850 12418 11159
rect 12670 11074 12698 11551
rect 13006 11578 13034 11583
rect 13230 11578 13258 11583
rect 13006 11577 13258 11578
rect 13006 11551 13007 11577
rect 13033 11551 13231 11577
rect 13257 11551 13258 11577
rect 13006 11550 13258 11551
rect 13006 11545 13034 11550
rect 13230 11545 13258 11550
rect 12726 11521 12754 11527
rect 12726 11495 12727 11521
rect 12753 11495 12754 11521
rect 12726 11241 12754 11495
rect 12726 11215 12727 11241
rect 12753 11215 12754 11241
rect 12726 11209 12754 11215
rect 13342 11242 13370 11607
rect 13342 11209 13370 11214
rect 13398 11577 13426 11583
rect 13398 11551 13399 11577
rect 13425 11551 13426 11577
rect 12670 11041 12698 11046
rect 13118 11074 13146 11079
rect 12390 10817 12418 10822
rect 12894 10850 12922 10855
rect 12110 10794 12138 10799
rect 12110 10747 12138 10766
rect 12614 10794 12642 10799
rect 12054 10430 12250 10458
rect 11886 9618 11914 9623
rect 11886 9571 11914 9590
rect 12166 9618 12194 9623
rect 12166 9571 12194 9590
rect 12110 9562 12138 9567
rect 12110 9515 12138 9534
rect 11774 9505 11802 9511
rect 11774 9479 11775 9505
rect 11801 9479 11802 9505
rect 11774 9450 11802 9479
rect 11774 9417 11802 9422
rect 11830 9505 11858 9511
rect 11830 9479 11831 9505
rect 11857 9479 11858 9505
rect 11830 9282 11858 9479
rect 11998 9506 12026 9511
rect 11998 9459 12026 9478
rect 11830 9249 11858 9254
rect 12166 9282 12194 9287
rect 11774 8721 11802 8727
rect 11774 8695 11775 8721
rect 11801 8695 11802 8721
rect 11774 8161 11802 8695
rect 11774 8135 11775 8161
rect 11801 8135 11802 8161
rect 11774 8129 11802 8135
rect 11886 8050 11914 8055
rect 10990 7713 11298 7714
rect 10990 7687 10991 7713
rect 11017 7687 11298 7713
rect 10990 7686 11298 7687
rect 10990 7681 11018 7686
rect 11270 7658 11298 7686
rect 11494 8049 11914 8050
rect 11494 8023 11887 8049
rect 11913 8023 11914 8049
rect 11494 8022 11914 8023
rect 11382 7658 11410 7663
rect 11270 7657 11410 7658
rect 11270 7631 11383 7657
rect 11409 7631 11410 7657
rect 11270 7630 11410 7631
rect 11382 7625 11410 7630
rect 11494 7657 11522 8022
rect 11886 8017 11914 8022
rect 11998 8049 12026 8055
rect 11998 8023 11999 8049
rect 12025 8023 12026 8049
rect 11494 7631 11495 7657
rect 11521 7631 11522 7657
rect 11494 7625 11522 7631
rect 11942 7937 11970 7943
rect 11942 7911 11943 7937
rect 11969 7911 11970 7937
rect 10822 7546 10906 7574
rect 11326 7546 11354 7551
rect 10766 7351 10767 7377
rect 10793 7351 10794 7377
rect 10766 7345 10794 7351
rect 10878 7378 10906 7546
rect 10878 7331 10906 7350
rect 11214 7545 11354 7546
rect 11214 7519 11327 7545
rect 11353 7519 11354 7545
rect 11214 7518 11354 7519
rect 10374 7321 10402 7327
rect 10374 7295 10375 7321
rect 10401 7295 10402 7321
rect 10374 7266 10402 7295
rect 10654 7266 10682 7271
rect 10374 7265 10682 7266
rect 10374 7239 10655 7265
rect 10681 7239 10682 7265
rect 10374 7238 10682 7239
rect 9534 7233 9562 7238
rect 10206 7219 10234 7238
rect 10654 7233 10682 7238
rect 9646 7154 9674 7159
rect 9646 6929 9674 7126
rect 9646 6903 9647 6929
rect 9673 6903 9674 6929
rect 9646 6897 9674 6903
rect 9814 7153 9842 7159
rect 9814 7127 9815 7153
rect 9841 7127 9842 7153
rect 9310 6827 9338 6846
rect 8974 6511 8975 6537
rect 9001 6511 9002 6537
rect 8974 6505 9002 6511
rect 9814 6370 9842 7127
rect 10318 7154 10346 7159
rect 10710 7154 10738 7159
rect 10318 7153 10402 7154
rect 10318 7127 10319 7153
rect 10345 7127 10402 7153
rect 10318 7126 10402 7127
rect 10318 7121 10346 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10318 6874 10346 6879
rect 10038 6537 10066 6543
rect 10038 6511 10039 6537
rect 10065 6511 10066 6537
rect 10038 6370 10066 6511
rect 10318 6537 10346 6846
rect 10374 6818 10402 7126
rect 10710 7107 10738 7126
rect 11214 6930 11242 7518
rect 11326 7513 11354 7518
rect 11550 7545 11578 7551
rect 11550 7519 11551 7545
rect 11577 7519 11578 7545
rect 11438 7378 11466 7383
rect 11550 7378 11578 7519
rect 11438 7377 11578 7378
rect 11438 7351 11439 7377
rect 11465 7351 11578 7377
rect 11438 7350 11578 7351
rect 11438 7345 11466 7350
rect 11942 7322 11970 7911
rect 11998 7882 12026 8023
rect 12166 7993 12194 9254
rect 12222 9226 12250 10430
rect 12614 10065 12642 10766
rect 12894 10793 12922 10822
rect 12894 10767 12895 10793
rect 12921 10767 12922 10793
rect 12894 10457 12922 10767
rect 12894 10431 12895 10457
rect 12921 10431 12922 10457
rect 12614 10039 12615 10065
rect 12641 10039 12642 10065
rect 12614 10033 12642 10039
rect 12782 10065 12810 10071
rect 12782 10039 12783 10065
rect 12809 10039 12810 10065
rect 12782 10010 12810 10039
rect 12782 9977 12810 9982
rect 12894 9617 12922 10431
rect 13118 10121 13146 11046
rect 13286 10738 13314 10743
rect 13118 10095 13119 10121
rect 13145 10095 13146 10121
rect 13118 10089 13146 10095
rect 13174 10737 13314 10738
rect 13174 10711 13287 10737
rect 13313 10711 13314 10737
rect 13174 10710 13314 10711
rect 13174 10121 13202 10710
rect 13286 10705 13314 10710
rect 13174 10095 13175 10121
rect 13201 10095 13202 10121
rect 13174 10089 13202 10095
rect 13398 10066 13426 11551
rect 13790 11242 13818 11247
rect 13790 11195 13818 11214
rect 14014 11241 14042 11998
rect 14294 12026 14322 12031
rect 14294 11979 14322 11998
rect 14574 12026 14602 12031
rect 14574 11969 14602 11998
rect 14686 11970 14714 12558
rect 15078 12026 15106 13063
rect 15302 13034 15330 13039
rect 15302 12305 15330 13006
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 18830 12698 18858 13119
rect 18942 13034 18970 13511
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 18942 13001 18970 13006
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 18830 12665 18858 12670
rect 15302 12279 15303 12305
rect 15329 12279 15330 12305
rect 15302 12273 15330 12279
rect 18830 12361 18858 12367
rect 18830 12335 18831 12361
rect 18857 12335 18858 12361
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 15078 11993 15106 11998
rect 15190 12026 15218 12031
rect 14574 11943 14575 11969
rect 14601 11943 14602 11969
rect 14574 11937 14602 11943
rect 14630 11942 14714 11970
rect 14630 11578 14658 11942
rect 14966 11914 14994 11919
rect 14686 11913 14994 11914
rect 14686 11887 14967 11913
rect 14993 11887 14994 11913
rect 14686 11886 14994 11887
rect 14686 11689 14714 11886
rect 14966 11881 14994 11886
rect 14686 11663 14687 11689
rect 14713 11663 14714 11689
rect 14686 11657 14714 11663
rect 14798 11690 14826 11695
rect 14798 11643 14826 11662
rect 15190 11689 15218 11998
rect 16030 12026 16058 12031
rect 16030 11979 16058 11998
rect 18830 12026 18858 12335
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 18830 11993 18858 11998
rect 15190 11663 15191 11689
rect 15217 11663 15218 11689
rect 15190 11657 15218 11663
rect 14686 11578 14714 11583
rect 14630 11550 14686 11578
rect 14014 11215 14015 11241
rect 14041 11215 14042 11241
rect 14014 10906 14042 11215
rect 14014 10873 14042 10878
rect 14630 10906 14658 10911
rect 14518 10793 14546 10799
rect 14518 10767 14519 10793
rect 14545 10767 14546 10793
rect 13398 10033 13426 10038
rect 14070 10738 14098 10743
rect 14070 10065 14098 10710
rect 14350 10738 14378 10743
rect 14350 10691 14378 10710
rect 14518 10094 14546 10767
rect 14070 10039 14071 10065
rect 14097 10039 14098 10065
rect 14070 10033 14098 10039
rect 14126 10066 14154 10071
rect 14126 10019 14154 10038
rect 14350 10065 14378 10071
rect 14350 10039 14351 10065
rect 14377 10039 14378 10065
rect 13230 10010 13258 10015
rect 13258 9982 13314 10010
rect 13230 9963 13258 9982
rect 13230 9674 13258 9679
rect 13230 9627 13258 9646
rect 12894 9591 12895 9617
rect 12921 9591 12922 9617
rect 12894 9585 12922 9591
rect 12838 9338 12866 9343
rect 12838 9291 12866 9310
rect 12222 8945 12250 9198
rect 12558 9282 12586 9287
rect 12222 8919 12223 8945
rect 12249 8919 12250 8945
rect 12222 8913 12250 8919
rect 12502 9002 12530 9007
rect 12334 8890 12362 8895
rect 12334 8843 12362 8862
rect 12502 8889 12530 8974
rect 12502 8863 12503 8889
rect 12529 8863 12530 8889
rect 12502 8857 12530 8863
rect 12558 8833 12586 9254
rect 12950 9282 12978 9287
rect 12950 9235 12978 9254
rect 12614 9226 12642 9231
rect 12614 9179 12642 9198
rect 13062 9226 13090 9231
rect 13062 9179 13090 9198
rect 13286 9225 13314 9982
rect 13454 10009 13482 10015
rect 13454 9983 13455 10009
rect 13481 9983 13482 10009
rect 13454 9954 13482 9983
rect 13454 9921 13482 9926
rect 13566 10009 13594 10015
rect 13566 9983 13567 10009
rect 13593 9983 13594 10009
rect 13566 9730 13594 9983
rect 13678 10010 13706 10015
rect 13678 9963 13706 9982
rect 13902 10010 13930 10015
rect 13902 9963 13930 9982
rect 13958 10009 13986 10015
rect 13958 9983 13959 10009
rect 13985 9983 13986 10009
rect 13566 9697 13594 9702
rect 13622 9953 13650 9959
rect 13622 9927 13623 9953
rect 13649 9927 13650 9953
rect 13622 9674 13650 9927
rect 13958 9954 13986 9983
rect 14238 10010 14266 10015
rect 14238 9963 14266 9982
rect 13958 9921 13986 9926
rect 13622 9641 13650 9646
rect 14294 9674 14322 9679
rect 14350 9674 14378 10039
rect 14406 10066 14546 10094
rect 14630 10401 14658 10878
rect 14630 10375 14631 10401
rect 14657 10375 14658 10401
rect 14406 10019 14434 10038
rect 14322 9646 14378 9674
rect 14630 9953 14658 10375
rect 14686 10849 14714 11550
rect 14854 11578 14882 11583
rect 15078 11578 15106 11583
rect 14854 11577 15106 11578
rect 14854 11551 14855 11577
rect 14881 11551 15079 11577
rect 15105 11551 15106 11577
rect 14854 11550 15106 11551
rect 14854 11545 14882 11550
rect 15078 11545 15106 11550
rect 15246 11578 15274 11583
rect 15246 11531 15274 11550
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 14910 10906 14938 10911
rect 14910 10859 14938 10878
rect 14686 10823 14687 10849
rect 14713 10823 14714 10849
rect 14686 10010 14714 10823
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10794 20034 10799
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 16086 10457 16114 10463
rect 16086 10431 16087 10457
rect 16113 10431 16114 10457
rect 16086 10402 16114 10431
rect 20006 10458 20034 10463
rect 20006 10411 20034 10430
rect 16310 10402 16338 10407
rect 16086 10401 16338 10402
rect 16086 10375 16311 10401
rect 16337 10375 16338 10401
rect 16086 10374 16338 10375
rect 15022 10346 15050 10351
rect 14854 10345 15050 10346
rect 14854 10319 15023 10345
rect 15049 10319 15050 10345
rect 14854 10318 15050 10319
rect 14854 10121 14882 10318
rect 15022 10313 15050 10318
rect 14854 10095 14855 10121
rect 14881 10095 14882 10121
rect 14854 10089 14882 10095
rect 14686 9977 14714 9982
rect 14966 10065 14994 10071
rect 14966 10039 14967 10065
rect 14993 10039 14994 10065
rect 14630 9927 14631 9953
rect 14657 9927 14658 9953
rect 14294 9627 14322 9646
rect 14630 9506 14658 9927
rect 14630 9505 14714 9506
rect 14630 9479 14631 9505
rect 14657 9479 14714 9505
rect 14630 9478 14714 9479
rect 14630 9473 14658 9478
rect 13286 9199 13287 9225
rect 13313 9199 13314 9225
rect 13118 9170 13146 9175
rect 13118 9123 13146 9142
rect 12670 9113 12698 9119
rect 12670 9087 12671 9113
rect 12697 9087 12698 9113
rect 12670 8946 12698 9087
rect 13286 9058 13314 9199
rect 12894 9030 13314 9058
rect 13398 9225 13426 9231
rect 13398 9199 13399 9225
rect 13425 9199 13426 9225
rect 13398 9114 13426 9199
rect 13454 9225 13482 9231
rect 13454 9199 13455 9225
rect 13481 9199 13482 9225
rect 13454 9170 13482 9199
rect 13454 9137 13482 9142
rect 12670 8913 12698 8918
rect 12782 9002 12810 9007
rect 12558 8807 12559 8833
rect 12585 8807 12586 8833
rect 12558 8801 12586 8807
rect 12782 8833 12810 8974
rect 12782 8807 12783 8833
rect 12809 8807 12810 8833
rect 12782 8801 12810 8807
rect 12894 8833 12922 9030
rect 12894 8807 12895 8833
rect 12921 8807 12922 8833
rect 12894 8801 12922 8807
rect 12950 8834 12978 8839
rect 12950 8787 12978 8806
rect 13398 8834 13426 9086
rect 13678 9114 13706 9119
rect 13678 9113 13818 9114
rect 13678 9087 13679 9113
rect 13705 9087 13818 9113
rect 13678 9086 13818 9087
rect 13678 9081 13706 9086
rect 13398 8801 13426 8806
rect 13790 8833 13818 9086
rect 13790 8807 13791 8833
rect 13817 8807 13818 8833
rect 13790 8801 13818 8807
rect 12446 8721 12474 8727
rect 12446 8695 12447 8721
rect 12473 8695 12474 8721
rect 12446 8162 12474 8695
rect 13174 8722 13202 8727
rect 13174 8721 13426 8722
rect 13174 8695 13175 8721
rect 13201 8695 13426 8721
rect 13174 8694 13426 8695
rect 13174 8689 13202 8694
rect 13398 8497 13426 8694
rect 13958 8721 13986 8727
rect 13958 8695 13959 8721
rect 13985 8695 13986 8721
rect 13398 8471 13399 8497
rect 13425 8471 13426 8497
rect 13398 8465 13426 8471
rect 13566 8497 13594 8503
rect 13566 8471 13567 8497
rect 13593 8471 13594 8497
rect 12446 8129 12474 8134
rect 12166 7967 12167 7993
rect 12193 7967 12194 7993
rect 12166 7961 12194 7967
rect 12222 7937 12250 7943
rect 12222 7911 12223 7937
rect 12249 7911 12250 7937
rect 12222 7882 12250 7911
rect 12278 7938 12306 7943
rect 12278 7891 12306 7910
rect 12782 7938 12810 7943
rect 11998 7854 12250 7882
rect 12782 7769 12810 7910
rect 12782 7743 12783 7769
rect 12809 7743 12810 7769
rect 12782 7602 12810 7743
rect 13286 7938 13314 7943
rect 12614 7546 12810 7574
rect 12950 7713 12978 7719
rect 12950 7687 12951 7713
rect 12977 7687 12978 7713
rect 11998 7322 12026 7327
rect 11942 7321 12026 7322
rect 11942 7295 11999 7321
rect 12025 7295 12026 7321
rect 11942 7294 12026 7295
rect 11998 7289 12026 7294
rect 11270 7266 11298 7271
rect 11270 7219 11298 7238
rect 11438 7265 11466 7271
rect 11438 7239 11439 7265
rect 11465 7239 11466 7265
rect 11270 6930 11298 6935
rect 11214 6929 11298 6930
rect 11214 6903 11271 6929
rect 11297 6903 11298 6929
rect 11214 6902 11298 6903
rect 11270 6897 11298 6902
rect 10766 6874 10794 6879
rect 10934 6874 10962 6879
rect 10794 6846 10850 6874
rect 10766 6841 10794 6846
rect 10710 6818 10738 6823
rect 10374 6817 10738 6818
rect 10374 6791 10711 6817
rect 10737 6791 10738 6817
rect 10374 6790 10738 6791
rect 10318 6511 10319 6537
rect 10345 6511 10346 6537
rect 10318 6505 10346 6511
rect 9814 6342 10066 6370
rect 9814 5082 9842 6342
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9814 5049 9842 5054
rect 10206 5082 10234 5087
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 8694 2143 8695 2169
rect 8721 2143 8722 2169
rect 8694 2137 8722 2143
rect 10206 2169 10234 5054
rect 10206 2143 10207 2169
rect 10233 2143 10234 2169
rect 10206 2137 10234 2143
rect 9254 2114 9282 2119
rect 9254 2067 9282 2086
rect 8638 1751 8639 1777
rect 8665 1751 8666 1777
rect 8638 1745 8666 1751
rect 10094 2058 10122 2063
rect 8414 1722 8442 1727
rect 8414 400 8442 1694
rect 9030 1722 9058 1727
rect 9030 1665 9058 1694
rect 9030 1639 9031 1665
rect 9057 1639 9058 1665
rect 9030 1633 9058 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10094 400 10122 2030
rect 10654 1778 10682 6790
rect 10710 6785 10738 6790
rect 10822 6537 10850 6846
rect 10934 6827 10962 6846
rect 11438 6818 11466 7239
rect 11606 7265 11634 7271
rect 11606 7239 11607 7265
rect 11633 7239 11634 7265
rect 11606 6874 11634 7239
rect 11606 6841 11634 6846
rect 11438 6785 11466 6790
rect 12278 6818 12306 6823
rect 12334 6818 12362 6823
rect 12306 6817 12362 6818
rect 12306 6791 12335 6817
rect 12361 6791 12362 6817
rect 12306 6790 12362 6791
rect 10822 6511 10823 6537
rect 10849 6511 10850 6537
rect 10822 6505 10850 6511
rect 10710 2058 10738 2063
rect 10710 2011 10738 2030
rect 10766 1834 10794 1839
rect 10710 1778 10738 1783
rect 10654 1777 10738 1778
rect 10654 1751 10711 1777
rect 10737 1751 10738 1777
rect 10654 1750 10738 1751
rect 10710 1745 10738 1750
rect 10766 400 10794 1806
rect 11214 1834 11242 1839
rect 11214 1787 11242 1806
rect 11774 1834 11802 1839
rect 11774 400 11802 1806
rect 12278 1777 12306 6790
rect 12334 6785 12362 6790
rect 12614 2169 12642 7546
rect 12670 6874 12698 6879
rect 12670 6827 12698 6846
rect 12950 4214 12978 7687
rect 13286 7658 13314 7910
rect 13566 7714 13594 8471
rect 13958 8498 13986 8695
rect 13958 8465 13986 8470
rect 14294 8498 14322 8503
rect 14294 8451 14322 8470
rect 13902 8441 13930 8447
rect 13902 8415 13903 8441
rect 13929 8415 13930 8441
rect 13734 7938 13762 7943
rect 13902 7938 13930 8415
rect 14574 8162 14602 8167
rect 14574 8115 14602 8134
rect 13762 7910 13930 7938
rect 14630 7993 14658 7999
rect 14630 7967 14631 7993
rect 14657 7967 14658 7993
rect 13734 7891 13762 7910
rect 13734 7714 13762 7719
rect 13566 7713 13762 7714
rect 13566 7687 13735 7713
rect 13761 7687 13762 7713
rect 13566 7686 13762 7687
rect 13734 7681 13762 7686
rect 13342 7658 13370 7663
rect 13286 7657 13370 7658
rect 13286 7631 13343 7657
rect 13369 7631 13370 7657
rect 13286 7630 13370 7631
rect 13062 7602 13090 7607
rect 13062 7321 13090 7574
rect 13062 7295 13063 7321
rect 13089 7295 13090 7321
rect 13062 7289 13090 7295
rect 13286 7153 13314 7630
rect 13342 7625 13370 7630
rect 14630 7602 14658 7967
rect 14686 7938 14714 9478
rect 14910 9226 14938 9231
rect 14910 8945 14938 9198
rect 14966 9114 14994 10039
rect 15246 10066 15274 10071
rect 15246 10019 15274 10038
rect 15022 10010 15050 10015
rect 15134 10010 15162 10015
rect 15022 10009 15162 10010
rect 15022 9983 15023 10009
rect 15049 9983 15135 10009
rect 15161 9983 15162 10009
rect 15022 9982 15162 9983
rect 15022 9977 15050 9982
rect 15134 9977 15162 9982
rect 15302 10010 15330 10015
rect 15302 9963 15330 9982
rect 16310 10010 16338 10374
rect 16422 10402 16450 10407
rect 16422 10345 16450 10374
rect 18830 10402 18858 10407
rect 18830 10355 18858 10374
rect 16422 10319 16423 10345
rect 16449 10319 16450 10345
rect 16422 10313 16450 10319
rect 20006 10066 20034 10071
rect 16310 9977 16338 9982
rect 18830 10010 18858 10015
rect 18830 9963 18858 9982
rect 20006 9953 20034 10038
rect 20006 9927 20007 9953
rect 20033 9927 20034 9953
rect 20006 9921 20034 9927
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9786 20034 9791
rect 20006 9729 20034 9758
rect 20006 9703 20007 9729
rect 20033 9703 20034 9729
rect 20006 9697 20034 9703
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 14966 9081 14994 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 14910 8919 14911 8945
rect 14937 8919 14938 8945
rect 14910 8913 14938 8919
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 14966 8834 14994 8839
rect 14966 8787 14994 8806
rect 15358 8834 15386 8839
rect 15358 8385 15386 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 15358 8359 15359 8385
rect 15385 8359 15386 8385
rect 15358 8353 15386 8359
rect 18830 8441 18858 8447
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 14686 7905 14714 7910
rect 15022 7938 15050 7943
rect 15022 7769 15050 7910
rect 15022 7743 15023 7769
rect 15049 7743 15050 7769
rect 15022 7737 15050 7743
rect 14798 7602 14826 7607
rect 14630 7574 14798 7602
rect 14798 7555 14826 7574
rect 18830 7602 18858 8415
rect 20006 8442 20034 8447
rect 20006 8385 20034 8414
rect 20006 8359 20007 8385
rect 20033 8359 20034 8385
rect 20006 8353 20034 8359
rect 18830 7569 18858 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13286 7127 13287 7153
rect 13313 7127 13314 7153
rect 13286 6874 13314 7127
rect 13286 6841 13314 6846
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 12894 4186 12978 4214
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 12838 2618 12866 2623
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12446 2058 12474 2063
rect 12446 400 12474 2030
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12838 1218 12866 2590
rect 12894 2561 12922 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 13398 2618 13426 2623
rect 13398 2571 13426 2590
rect 12894 2535 12895 2561
rect 12921 2535 12922 2561
rect 12894 2529 12922 2535
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1190 12866 1218
rect 12782 400 12810 1190
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 10080 0 10136 400
rect 10752 0 10808 400
rect 11760 0 11816 400
rect 12432 0 12488 400
rect 12768 0 12824 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8414 19110 8442 19138
rect 9030 19137 9058 19138
rect 9030 19111 9031 19137
rect 9031 19111 9057 19137
rect 9057 19111 9058 19137
rect 9030 19110 9058 19111
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 10430 19110 10458 19138
rect 11046 19137 11074 19138
rect 11046 19111 11047 19137
rect 11047 19111 11073 19137
rect 11073 19111 11074 19137
rect 11046 19110 11074 19111
rect 12782 19278 12810 19306
rect 12110 19110 12138 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 13118 19110 13146 19138
rect 13398 19278 13426 19306
rect 10094 18718 10122 18746
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 2142 13537 2170 13538
rect 2142 13511 2143 13537
rect 2143 13511 2169 13537
rect 2169 13511 2170 13537
rect 2142 13510 2170 13511
rect 6062 13510 6090 13538
rect 966 13118 994 13146
rect 2086 13454 2114 13482
rect 966 12446 994 12474
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 7462 13398 7490 13426
rect 7854 13398 7882 13426
rect 7070 13174 7098 13202
rect 7406 13174 7434 13202
rect 8750 13174 8778 13202
rect 6062 13089 6090 13090
rect 6062 13063 6063 13089
rect 6063 13063 6089 13089
rect 6089 13063 6090 13089
rect 6062 13062 6090 13063
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 6958 12697 6986 12698
rect 6958 12671 6959 12697
rect 6959 12671 6985 12697
rect 6985 12671 6986 12697
rect 6958 12670 6986 12671
rect 7574 13062 7602 13090
rect 7518 12697 7546 12698
rect 7518 12671 7519 12697
rect 7519 12671 7545 12697
rect 7545 12671 7546 12697
rect 7518 12670 7546 12671
rect 7630 12697 7658 12698
rect 7630 12671 7631 12697
rect 7631 12671 7657 12697
rect 7657 12671 7658 12697
rect 7630 12670 7658 12671
rect 7406 12614 7434 12642
rect 6678 12446 6706 12474
rect 7686 12558 7714 12586
rect 7350 12473 7378 12474
rect 7350 12447 7351 12473
rect 7351 12447 7377 12473
rect 7377 12447 7378 12473
rect 7350 12446 7378 12447
rect 7294 12361 7322 12362
rect 7294 12335 7295 12361
rect 7295 12335 7321 12361
rect 7321 12335 7322 12361
rect 7294 12334 7322 12335
rect 2142 12278 2170 12306
rect 5614 12305 5642 12306
rect 5614 12279 5615 12305
rect 5615 12279 5641 12305
rect 5641 12279 5642 12305
rect 5614 12278 5642 12279
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 5614 11998 5642 12026
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 8078 12641 8106 12642
rect 8078 12615 8079 12641
rect 8079 12615 8105 12641
rect 8105 12615 8106 12641
rect 8078 12614 8106 12615
rect 7854 12446 7882 12474
rect 7126 12025 7154 12026
rect 7126 11999 7127 12025
rect 7127 11999 7153 12025
rect 7153 11999 7154 12025
rect 7126 11998 7154 11999
rect 7686 11662 7714 11690
rect 8302 12558 8330 12586
rect 8750 12614 8778 12642
rect 8022 12334 8050 12362
rect 7910 11662 7938 11690
rect 5614 11521 5642 11522
rect 5614 11495 5615 11521
rect 5615 11495 5641 11521
rect 5641 11495 5642 11521
rect 5614 11494 5642 11495
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6678 11521 6706 11522
rect 6678 11495 6679 11521
rect 6679 11495 6705 11521
rect 6705 11495 6706 11521
rect 6678 11494 6706 11495
rect 5614 11102 5642 11130
rect 6062 11046 6090 11074
rect 7406 11521 7434 11522
rect 7406 11495 7407 11521
rect 7407 11495 7433 11521
rect 7433 11495 7434 11521
rect 7406 11494 7434 11495
rect 7238 11185 7266 11186
rect 7238 11159 7239 11185
rect 7239 11159 7265 11185
rect 7265 11159 7266 11185
rect 7238 11158 7266 11159
rect 7182 11129 7210 11130
rect 7182 11103 7183 11129
rect 7183 11103 7209 11129
rect 7209 11103 7210 11129
rect 7182 11102 7210 11103
rect 7630 11270 7658 11298
rect 7798 11158 7826 11186
rect 7854 11214 7882 11242
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 7126 10737 7154 10738
rect 7126 10711 7127 10737
rect 7127 10711 7153 10737
rect 7153 10711 7154 10737
rect 7126 10710 7154 10711
rect 7350 10822 7378 10850
rect 5670 10094 5698 10122
rect 7462 10710 7490 10738
rect 7518 10513 7546 10514
rect 7518 10487 7519 10513
rect 7519 10487 7545 10513
rect 7545 10487 7546 10513
rect 7518 10486 7546 10487
rect 7686 11073 7714 11074
rect 7686 11047 7687 11073
rect 7687 11047 7713 11073
rect 7713 11047 7714 11073
rect 7686 11046 7714 11047
rect 7742 10486 7770 10514
rect 7238 10094 7266 10122
rect 7686 10094 7714 10122
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 2086 9478 2114 9506
rect 5950 9281 5978 9282
rect 5950 9255 5951 9281
rect 5951 9255 5977 9281
rect 5977 9255 5978 9281
rect 5950 9254 5978 9255
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 7350 10065 7378 10066
rect 7350 10039 7351 10065
rect 7351 10039 7377 10065
rect 7377 10039 7378 10065
rect 7350 10038 7378 10039
rect 7238 9310 7266 9338
rect 7014 9169 7042 9170
rect 7014 9143 7015 9169
rect 7015 9143 7041 9169
rect 7041 9143 7042 9169
rect 7014 9142 7042 9143
rect 6006 8750 6034 8778
rect 6902 8777 6930 8778
rect 6902 8751 6903 8777
rect 6903 8751 6929 8777
rect 6929 8751 6930 8777
rect 6902 8750 6930 8751
rect 7406 9310 7434 9338
rect 7630 10009 7658 10010
rect 7630 9983 7631 10009
rect 7631 9983 7657 10009
rect 7657 9983 7658 10009
rect 7630 9982 7658 9983
rect 7742 9870 7770 9898
rect 8638 12558 8666 12586
rect 8470 12502 8498 12530
rect 9030 12502 9058 12530
rect 8862 12361 8890 12362
rect 8862 12335 8863 12361
rect 8863 12335 8889 12361
rect 8889 12335 8890 12361
rect 8862 12334 8890 12335
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9310 12838 9338 12866
rect 10710 18745 10738 18746
rect 10710 18719 10711 18745
rect 10711 18719 10737 18745
rect 10737 18719 10738 18745
rect 10710 18718 10738 18719
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 14686 19137 14714 19138
rect 14686 19111 14687 19137
rect 14687 19111 14713 19137
rect 14713 19111 14714 19137
rect 14686 19110 14714 19111
rect 9702 12753 9730 12754
rect 9702 12727 9703 12753
rect 9703 12727 9729 12753
rect 9729 12727 9730 12753
rect 9702 12726 9730 12727
rect 9142 12446 9170 12474
rect 9198 12670 9226 12698
rect 8806 11942 8834 11970
rect 8526 11857 8554 11858
rect 8526 11831 8527 11857
rect 8527 11831 8553 11857
rect 8553 11831 8554 11857
rect 8526 11830 8554 11831
rect 9086 11886 9114 11914
rect 8918 11718 8946 11746
rect 8862 11689 8890 11690
rect 8862 11663 8863 11689
rect 8863 11663 8889 11689
rect 8889 11663 8890 11689
rect 8862 11662 8890 11663
rect 8022 11214 8050 11242
rect 7966 11158 7994 11186
rect 8358 10878 8386 10906
rect 8134 10542 8162 10570
rect 8078 10121 8106 10122
rect 8078 10095 8079 10121
rect 8079 10095 8105 10121
rect 8105 10095 8106 10121
rect 8078 10094 8106 10095
rect 8134 10038 8162 10066
rect 7910 9646 7938 9674
rect 8246 10038 8274 10066
rect 8750 10822 8778 10850
rect 8526 10401 8554 10402
rect 8526 10375 8527 10401
rect 8527 10375 8553 10401
rect 8553 10375 8554 10401
rect 8526 10374 8554 10375
rect 8302 9982 8330 10010
rect 7910 9561 7938 9562
rect 7910 9535 7911 9561
rect 7911 9535 7937 9561
rect 7937 9535 7938 9561
rect 7910 9534 7938 9535
rect 7742 9310 7770 9338
rect 8078 9254 8106 9282
rect 7350 9142 7378 9170
rect 8246 9142 8274 9170
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 8638 9982 8666 10010
rect 8974 11633 9002 11634
rect 8974 11607 8975 11633
rect 8975 11607 9001 11633
rect 9001 11607 9002 11633
rect 8974 11606 9002 11607
rect 9030 11214 9058 11242
rect 9086 10374 9114 10402
rect 9534 12502 9562 12530
rect 9758 12614 9786 12642
rect 9254 12390 9282 12418
rect 9254 11969 9282 11970
rect 9254 11943 9255 11969
rect 9255 11943 9281 11969
rect 9281 11943 9282 11969
rect 9254 11942 9282 11943
rect 10150 12782 10178 12810
rect 9870 12670 9898 12698
rect 9982 12697 10010 12698
rect 9982 12671 9983 12697
rect 9983 12671 10009 12697
rect 10009 12671 10010 12697
rect 9982 12670 10010 12671
rect 10094 12614 10122 12642
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9814 12390 9842 12418
rect 9814 12249 9842 12250
rect 9814 12223 9815 12249
rect 9815 12223 9841 12249
rect 9841 12223 9842 12249
rect 9814 12222 9842 12223
rect 10318 13174 10346 13202
rect 10878 13174 10906 13202
rect 10710 13145 10738 13146
rect 10710 13119 10711 13145
rect 10711 13119 10737 13145
rect 10737 13119 10738 13145
rect 10710 13118 10738 13119
rect 10710 12838 10738 12866
rect 11774 13118 11802 13146
rect 12110 13230 12138 13258
rect 12334 13454 12362 13482
rect 13398 13481 13426 13482
rect 13398 13455 13399 13481
rect 13399 13455 13425 13481
rect 13425 13455 13426 13481
rect 13398 13454 13426 13455
rect 12670 13257 12698 13258
rect 12670 13231 12671 13257
rect 12671 13231 12697 13257
rect 12697 13231 12698 13257
rect 12670 13230 12698 13231
rect 12726 13201 12754 13202
rect 12726 13175 12727 13201
rect 12727 13175 12753 13201
rect 12753 13175 12754 13201
rect 12726 13174 12754 13175
rect 13118 13257 13146 13258
rect 13118 13231 13119 13257
rect 13119 13231 13145 13257
rect 13145 13231 13146 13257
rect 13118 13230 13146 13231
rect 12334 13145 12362 13146
rect 12334 13119 12335 13145
rect 12335 13119 12361 13145
rect 12361 13119 12362 13145
rect 12334 13118 12362 13119
rect 10822 12782 10850 12810
rect 10206 12726 10234 12754
rect 10654 12697 10682 12698
rect 10654 12671 10655 12697
rect 10655 12671 10681 12697
rect 10681 12671 10682 12697
rect 10654 12670 10682 12671
rect 10766 12641 10794 12642
rect 10766 12615 10767 12641
rect 10767 12615 10793 12641
rect 10793 12615 10794 12641
rect 10766 12614 10794 12615
rect 10206 12446 10234 12474
rect 10486 12222 10514 12250
rect 10430 12054 10458 12082
rect 9534 11886 9562 11914
rect 9590 11830 9618 11858
rect 9534 11633 9562 11634
rect 9534 11607 9535 11633
rect 9535 11607 9561 11633
rect 9561 11607 9562 11633
rect 9534 11606 9562 11607
rect 9534 11214 9562 11242
rect 9310 10878 9338 10906
rect 9254 10849 9282 10850
rect 9254 10823 9255 10849
rect 9255 10823 9281 10849
rect 9281 10823 9282 10849
rect 9254 10822 9282 10823
rect 9254 10542 9282 10570
rect 9870 11913 9898 11914
rect 9870 11887 9871 11913
rect 9871 11887 9897 11913
rect 9897 11887 9898 11913
rect 9870 11886 9898 11887
rect 9814 11830 9842 11858
rect 9982 11857 10010 11858
rect 9982 11831 9983 11857
rect 9983 11831 10009 11857
rect 10009 11831 10010 11857
rect 9982 11830 10010 11831
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10094 11718 10122 11746
rect 9758 11521 9786 11522
rect 9758 11495 9759 11521
rect 9759 11495 9785 11521
rect 9785 11495 9786 11521
rect 9758 11494 9786 11495
rect 9534 11046 9562 11074
rect 8806 9870 8834 9898
rect 8918 10009 8946 10010
rect 8918 9983 8919 10009
rect 8919 9983 8945 10009
rect 8945 9983 8946 10009
rect 8918 9982 8946 9983
rect 8862 9729 8890 9730
rect 8862 9703 8863 9729
rect 8863 9703 8889 9729
rect 8889 9703 8890 9729
rect 8862 9702 8890 9703
rect 8862 9590 8890 9618
rect 8806 9561 8834 9562
rect 8806 9535 8807 9561
rect 8807 9535 8833 9561
rect 8833 9535 8834 9561
rect 8806 9534 8834 9535
rect 8974 9953 9002 9954
rect 8974 9927 8975 9953
rect 8975 9927 9001 9953
rect 9001 9927 9002 9953
rect 8974 9926 9002 9927
rect 9198 10094 9226 10122
rect 9366 9982 9394 10010
rect 9310 9926 9338 9954
rect 9142 9590 9170 9618
rect 8862 9254 8890 9282
rect 9030 9422 9058 9450
rect 8806 8833 8834 8834
rect 8806 8807 8807 8833
rect 8807 8807 8833 8833
rect 8833 8807 8834 8833
rect 8806 8806 8834 8807
rect 8974 8414 9002 8442
rect 8302 7910 8330 7938
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8414 7937 8442 7938
rect 8414 7911 8415 7937
rect 8415 7911 8441 7937
rect 8441 7911 8442 7937
rect 8414 7910 8442 7911
rect 9422 9953 9450 9954
rect 9422 9927 9423 9953
rect 9423 9927 9449 9953
rect 9449 9927 9450 9953
rect 9422 9926 9450 9927
rect 9422 9086 9450 9114
rect 9702 11185 9730 11186
rect 9702 11159 9703 11185
rect 9703 11159 9729 11185
rect 9729 11159 9730 11185
rect 9702 11158 9730 11159
rect 9646 10878 9674 10906
rect 9982 11046 10010 11074
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10262 11494 10290 11522
rect 9814 10542 9842 10570
rect 10374 11158 10402 11186
rect 10150 10542 10178 10570
rect 10542 11550 10570 11578
rect 11830 12726 11858 12754
rect 11102 12614 11130 12642
rect 11550 12697 11578 12698
rect 11550 12671 11551 12697
rect 11551 12671 11577 12697
rect 11577 12671 11578 12697
rect 11550 12670 11578 12671
rect 11494 12054 11522 12082
rect 11774 12614 11802 12642
rect 10766 11886 10794 11914
rect 10654 11718 10682 11746
rect 10542 11158 10570 11186
rect 10598 11270 10626 11298
rect 10710 11494 10738 11522
rect 10822 11857 10850 11858
rect 10822 11831 10823 11857
rect 10823 11831 10849 11857
rect 10849 11831 10850 11857
rect 10822 11830 10850 11831
rect 10598 10822 10626 10850
rect 9870 10289 9898 10290
rect 9870 10263 9871 10289
rect 9871 10263 9897 10289
rect 9897 10263 9898 10289
rect 9870 10262 9898 10263
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9758 10038 9786 10066
rect 10374 9982 10402 10010
rect 9758 9590 9786 9618
rect 9590 9478 9618 9506
rect 9590 9169 9618 9170
rect 9590 9143 9591 9169
rect 9591 9143 9617 9169
rect 9617 9143 9618 9169
rect 9590 9142 9618 9143
rect 9758 9198 9786 9226
rect 9702 9142 9730 9170
rect 9478 8750 9506 8778
rect 10206 9617 10234 9618
rect 10206 9591 10207 9617
rect 10207 9591 10233 9617
rect 10233 9591 10234 9617
rect 10206 9590 10234 9591
rect 9926 9561 9954 9562
rect 9926 9535 9927 9561
rect 9927 9535 9953 9561
rect 9953 9535 9954 9561
rect 9926 9534 9954 9535
rect 10038 9478 10066 9506
rect 10150 9534 10178 9562
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9870 9225 9898 9226
rect 9870 9199 9871 9225
rect 9871 9199 9897 9225
rect 9897 9199 9898 9225
rect 9870 9198 9898 9199
rect 10206 9169 10234 9170
rect 10206 9143 10207 9169
rect 10207 9143 10233 9169
rect 10233 9143 10234 9169
rect 10206 9142 10234 9143
rect 11158 11942 11186 11970
rect 11158 11857 11186 11858
rect 11158 11831 11159 11857
rect 11159 11831 11185 11857
rect 11185 11831 11186 11857
rect 11158 11830 11186 11831
rect 10990 11577 11018 11578
rect 10990 11551 10991 11577
rect 10991 11551 11017 11577
rect 11017 11551 11018 11577
rect 10990 11550 11018 11551
rect 10822 11102 10850 11130
rect 10766 10822 10794 10850
rect 10990 11129 11018 11130
rect 10990 11103 10991 11129
rect 10991 11103 11017 11129
rect 11017 11103 11018 11129
rect 10990 11102 11018 11103
rect 11326 11718 11354 11746
rect 11494 11606 11522 11634
rect 12334 12753 12362 12754
rect 12334 12727 12335 12753
rect 12335 12727 12361 12753
rect 12361 12727 12362 12753
rect 12334 12726 12362 12727
rect 12110 12670 12138 12698
rect 12390 12697 12418 12698
rect 12390 12671 12391 12697
rect 12391 12671 12417 12697
rect 12417 12671 12418 12697
rect 12390 12670 12418 12671
rect 12278 12614 12306 12642
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 14294 13230 14322 13258
rect 12950 12697 12978 12698
rect 12950 12671 12951 12697
rect 12951 12671 12977 12697
rect 12977 12671 12978 12697
rect 12950 12670 12978 12671
rect 14238 12726 14266 12754
rect 13790 12697 13818 12698
rect 13790 12671 13791 12697
rect 13791 12671 13817 12697
rect 13817 12671 13818 12697
rect 13790 12670 13818 12671
rect 14518 12697 14546 12698
rect 14518 12671 14519 12697
rect 14519 12671 14545 12697
rect 14545 12671 14546 12697
rect 14518 12670 14546 12671
rect 14630 12697 14658 12698
rect 14630 12671 14631 12697
rect 14631 12671 14657 12697
rect 14657 12671 14658 12697
rect 14630 12670 14658 12671
rect 13734 12641 13762 12642
rect 13734 12615 13735 12641
rect 13735 12615 13761 12641
rect 13761 12615 13762 12641
rect 13734 12614 13762 12615
rect 12782 12278 12810 12306
rect 14854 12670 14882 12698
rect 14910 13006 14938 13034
rect 13846 11998 13874 12026
rect 14014 11998 14042 12026
rect 11830 11633 11858 11634
rect 11830 11607 11831 11633
rect 11831 11607 11857 11633
rect 11857 11607 11858 11633
rect 11830 11606 11858 11607
rect 11494 11129 11522 11130
rect 11494 11103 11495 11129
rect 11495 11103 11521 11129
rect 11521 11103 11522 11129
rect 11494 11102 11522 11103
rect 11270 10878 11298 10906
rect 11214 10486 11242 10514
rect 10598 9926 10626 9954
rect 10710 10318 10738 10346
rect 10598 9310 10626 9338
rect 10654 9142 10682 9170
rect 10710 8833 10738 8834
rect 10710 8807 10711 8833
rect 10711 8807 10737 8833
rect 10737 8807 10738 8833
rect 10710 8806 10738 8807
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9814 8441 9842 8442
rect 9814 8415 9815 8441
rect 9815 8415 9841 8441
rect 9841 8415 9842 8441
rect 9814 8414 9842 8415
rect 9926 8497 9954 8498
rect 9926 8471 9927 8497
rect 9927 8471 9953 8497
rect 9953 8471 9954 8497
rect 9926 8470 9954 8471
rect 8694 7937 8722 7938
rect 8694 7911 8695 7937
rect 8695 7911 8721 7937
rect 8721 7911 8722 7937
rect 8694 7910 8722 7911
rect 9254 7910 9282 7938
rect 8302 7630 8330 7658
rect 7182 7574 7210 7602
rect 7238 7350 7266 7378
rect 8638 7630 8666 7658
rect 8470 7350 8498 7378
rect 8246 7321 8274 7322
rect 8246 7295 8247 7321
rect 8247 7295 8273 7321
rect 8273 7295 8274 7321
rect 8246 7294 8274 7295
rect 8582 7350 8610 7378
rect 6902 7238 6930 7266
rect 8358 7238 8386 7266
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8078 2086 8106 2114
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 8750 7601 8778 7602
rect 8750 7575 8751 7601
rect 8751 7575 8777 7601
rect 8777 7575 8778 7601
rect 8750 7574 8778 7575
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 8974 7350 9002 7378
rect 9310 7377 9338 7378
rect 9310 7351 9311 7377
rect 9311 7351 9337 7377
rect 9337 7351 9338 7377
rect 9310 7350 9338 7351
rect 8694 7294 8722 7322
rect 9086 7294 9114 7322
rect 8806 7265 8834 7266
rect 8806 7239 8807 7265
rect 8807 7239 8833 7265
rect 8833 7239 8834 7265
rect 8806 7238 8834 7239
rect 9310 7238 9338 7266
rect 8974 7182 9002 7210
rect 9254 7209 9282 7210
rect 9254 7183 9255 7209
rect 9255 7183 9281 7209
rect 9281 7183 9282 7209
rect 9254 7182 9282 7183
rect 10878 10318 10906 10346
rect 10822 10038 10850 10066
rect 10878 9590 10906 9618
rect 10934 9478 10962 9506
rect 10990 9225 11018 9226
rect 10990 9199 10991 9225
rect 10991 9199 11017 9225
rect 11017 9199 11018 9225
rect 10990 9198 11018 9199
rect 11326 10374 11354 10402
rect 11102 10262 11130 10290
rect 11158 9982 11186 10010
rect 11214 9534 11242 9562
rect 11326 8862 11354 8890
rect 11662 10793 11690 10794
rect 11662 10767 11663 10793
rect 11663 10767 11689 10793
rect 11689 10767 11690 10793
rect 11662 10766 11690 10767
rect 11550 10486 11578 10514
rect 11494 10038 11522 10066
rect 11662 10401 11690 10402
rect 11662 10375 11663 10401
rect 11663 10375 11689 10401
rect 11689 10375 11690 10401
rect 11662 10374 11690 10375
rect 11550 9870 11578 9898
rect 11550 9422 11578 9450
rect 11662 9478 11690 9506
rect 11494 9086 11522 9114
rect 11494 8806 11522 8834
rect 11046 8470 11074 8498
rect 12054 11550 12082 11578
rect 11998 11214 12026 11242
rect 11942 10905 11970 10906
rect 11942 10879 11943 10905
rect 11943 10879 11969 10905
rect 11969 10879 11970 10905
rect 11942 10878 11970 10879
rect 12166 11073 12194 11074
rect 12166 11047 12167 11073
rect 12167 11047 12193 11073
rect 12193 11047 12194 11073
rect 12166 11046 12194 11047
rect 13342 11214 13370 11242
rect 12670 11046 12698 11074
rect 13118 11046 13146 11074
rect 12390 10822 12418 10850
rect 12894 10822 12922 10850
rect 12110 10793 12138 10794
rect 12110 10767 12111 10793
rect 12111 10767 12137 10793
rect 12137 10767 12138 10793
rect 12110 10766 12138 10767
rect 12614 10766 12642 10794
rect 11886 9617 11914 9618
rect 11886 9591 11887 9617
rect 11887 9591 11913 9617
rect 11913 9591 11914 9617
rect 11886 9590 11914 9591
rect 12166 9617 12194 9618
rect 12166 9591 12167 9617
rect 12167 9591 12193 9617
rect 12193 9591 12194 9617
rect 12166 9590 12194 9591
rect 12110 9561 12138 9562
rect 12110 9535 12111 9561
rect 12111 9535 12137 9561
rect 12137 9535 12138 9561
rect 12110 9534 12138 9535
rect 11774 9422 11802 9450
rect 11998 9505 12026 9506
rect 11998 9479 11999 9505
rect 11999 9479 12025 9505
rect 12025 9479 12026 9505
rect 11998 9478 12026 9479
rect 11830 9254 11858 9282
rect 12166 9254 12194 9282
rect 10878 7377 10906 7378
rect 10878 7351 10879 7377
rect 10879 7351 10905 7377
rect 10905 7351 10906 7377
rect 10878 7350 10906 7351
rect 10206 7265 10234 7266
rect 10206 7239 10207 7265
rect 10207 7239 10233 7265
rect 10233 7239 10234 7265
rect 10206 7238 10234 7239
rect 9646 7126 9674 7154
rect 9310 6873 9338 6874
rect 9310 6847 9311 6873
rect 9311 6847 9337 6873
rect 9337 6847 9338 6873
rect 9310 6846 9338 6847
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10318 6846 10346 6874
rect 10710 7153 10738 7154
rect 10710 7127 10711 7153
rect 10711 7127 10737 7153
rect 10737 7127 10738 7153
rect 10710 7126 10738 7127
rect 12782 9982 12810 10010
rect 13790 11241 13818 11242
rect 13790 11215 13791 11241
rect 13791 11215 13817 11241
rect 13817 11215 13818 11241
rect 13790 11214 13818 11215
rect 14294 12025 14322 12026
rect 14294 11999 14295 12025
rect 14295 11999 14321 12025
rect 14321 11999 14322 12025
rect 14294 11998 14322 11999
rect 14574 11998 14602 12026
rect 15302 13006 15330 13034
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 20006 13118 20034 13146
rect 18942 13006 18970 13034
rect 20006 12782 20034 12810
rect 18830 12670 18858 12698
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 15078 11998 15106 12026
rect 15190 11998 15218 12026
rect 14798 11689 14826 11690
rect 14798 11663 14799 11689
rect 14799 11663 14825 11689
rect 14825 11663 14826 11689
rect 14798 11662 14826 11663
rect 16030 12025 16058 12026
rect 16030 11999 16031 12025
rect 16031 11999 16057 12025
rect 16057 11999 16058 12025
rect 16030 11998 16058 11999
rect 20006 12110 20034 12138
rect 18830 11998 18858 12026
rect 14686 11550 14714 11578
rect 14014 10878 14042 10906
rect 14630 10878 14658 10906
rect 13398 10038 13426 10066
rect 14070 10710 14098 10738
rect 14350 10737 14378 10738
rect 14350 10711 14351 10737
rect 14351 10711 14377 10737
rect 14377 10711 14378 10737
rect 14350 10710 14378 10711
rect 14126 10065 14154 10066
rect 14126 10039 14127 10065
rect 14127 10039 14153 10065
rect 14153 10039 14154 10065
rect 14126 10038 14154 10039
rect 13230 10009 13258 10010
rect 13230 9983 13231 10009
rect 13231 9983 13257 10009
rect 13257 9983 13258 10009
rect 13230 9982 13258 9983
rect 13230 9673 13258 9674
rect 13230 9647 13231 9673
rect 13231 9647 13257 9673
rect 13257 9647 13258 9673
rect 13230 9646 13258 9647
rect 12838 9337 12866 9338
rect 12838 9311 12839 9337
rect 12839 9311 12865 9337
rect 12865 9311 12866 9337
rect 12838 9310 12866 9311
rect 12222 9198 12250 9226
rect 12558 9254 12586 9282
rect 12502 8974 12530 9002
rect 12334 8889 12362 8890
rect 12334 8863 12335 8889
rect 12335 8863 12361 8889
rect 12361 8863 12362 8889
rect 12334 8862 12362 8863
rect 12950 9281 12978 9282
rect 12950 9255 12951 9281
rect 12951 9255 12977 9281
rect 12977 9255 12978 9281
rect 12950 9254 12978 9255
rect 12614 9225 12642 9226
rect 12614 9199 12615 9225
rect 12615 9199 12641 9225
rect 12641 9199 12642 9225
rect 12614 9198 12642 9199
rect 13062 9225 13090 9226
rect 13062 9199 13063 9225
rect 13063 9199 13089 9225
rect 13089 9199 13090 9225
rect 13062 9198 13090 9199
rect 13454 9926 13482 9954
rect 13678 10009 13706 10010
rect 13678 9983 13679 10009
rect 13679 9983 13705 10009
rect 13705 9983 13706 10009
rect 13678 9982 13706 9983
rect 13902 10009 13930 10010
rect 13902 9983 13903 10009
rect 13903 9983 13929 10009
rect 13929 9983 13930 10009
rect 13902 9982 13930 9983
rect 13566 9702 13594 9730
rect 14238 10009 14266 10010
rect 14238 9983 14239 10009
rect 14239 9983 14265 10009
rect 14265 9983 14266 10009
rect 14238 9982 14266 9983
rect 13958 9926 13986 9954
rect 13622 9646 13650 9674
rect 14406 10065 14434 10066
rect 14406 10039 14407 10065
rect 14407 10039 14433 10065
rect 14433 10039 14434 10065
rect 14406 10038 14434 10039
rect 14294 9673 14322 9674
rect 14294 9647 14295 9673
rect 14295 9647 14321 9673
rect 14321 9647 14322 9673
rect 14294 9646 14322 9647
rect 15246 11577 15274 11578
rect 15246 11551 15247 11577
rect 15247 11551 15273 11577
rect 15273 11551 15274 11577
rect 15246 11550 15274 11551
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 20006 11102 20034 11130
rect 14910 10905 14938 10906
rect 14910 10879 14911 10905
rect 14911 10879 14937 10905
rect 14937 10879 14938 10905
rect 14910 10878 14938 10879
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20006 10766 20034 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 20006 10457 20034 10458
rect 20006 10431 20007 10457
rect 20007 10431 20033 10457
rect 20033 10431 20034 10457
rect 20006 10430 20034 10431
rect 14686 9982 14714 10010
rect 13118 9169 13146 9170
rect 13118 9143 13119 9169
rect 13119 9143 13145 9169
rect 13145 9143 13146 9169
rect 13118 9142 13146 9143
rect 13454 9142 13482 9170
rect 13398 9086 13426 9114
rect 12670 8918 12698 8946
rect 12782 8974 12810 9002
rect 12950 8833 12978 8834
rect 12950 8807 12951 8833
rect 12951 8807 12977 8833
rect 12977 8807 12978 8833
rect 12950 8806 12978 8807
rect 13398 8806 13426 8834
rect 12446 8134 12474 8162
rect 12278 7937 12306 7938
rect 12278 7911 12279 7937
rect 12279 7911 12305 7937
rect 12305 7911 12306 7937
rect 12278 7910 12306 7911
rect 12782 7910 12810 7938
rect 13286 7910 13314 7938
rect 12782 7574 12810 7602
rect 11270 7265 11298 7266
rect 11270 7239 11271 7265
rect 11271 7239 11297 7265
rect 11297 7239 11298 7265
rect 11270 7238 11298 7239
rect 10766 6846 10794 6874
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9814 5054 9842 5082
rect 10206 5054 10234 5082
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9254 2113 9282 2114
rect 9254 2087 9255 2113
rect 9255 2087 9281 2113
rect 9281 2087 9282 2113
rect 9254 2086 9282 2087
rect 10094 2030 10122 2058
rect 8414 1694 8442 1722
rect 9030 1694 9058 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 10934 6873 10962 6874
rect 10934 6847 10935 6873
rect 10935 6847 10961 6873
rect 10961 6847 10962 6873
rect 10934 6846 10962 6847
rect 11606 6846 11634 6874
rect 11438 6790 11466 6818
rect 12278 6790 12306 6818
rect 10710 2057 10738 2058
rect 10710 2031 10711 2057
rect 10711 2031 10737 2057
rect 10737 2031 10738 2057
rect 10710 2030 10738 2031
rect 10766 1806 10794 1834
rect 11214 1833 11242 1834
rect 11214 1807 11215 1833
rect 11215 1807 11241 1833
rect 11241 1807 11242 1833
rect 11214 1806 11242 1807
rect 11774 1806 11802 1834
rect 12670 6873 12698 6874
rect 12670 6847 12671 6873
rect 12671 6847 12697 6873
rect 12697 6847 12698 6873
rect 12670 6846 12698 6847
rect 13958 8470 13986 8498
rect 14294 8497 14322 8498
rect 14294 8471 14295 8497
rect 14295 8471 14321 8497
rect 14321 8471 14322 8497
rect 14294 8470 14322 8471
rect 14574 8161 14602 8162
rect 14574 8135 14575 8161
rect 14575 8135 14601 8161
rect 14601 8135 14602 8161
rect 14574 8134 14602 8135
rect 13734 7937 13762 7938
rect 13734 7911 13735 7937
rect 13735 7911 13761 7937
rect 13761 7911 13762 7937
rect 13734 7910 13762 7911
rect 13062 7574 13090 7602
rect 14910 9198 14938 9226
rect 15246 10065 15274 10066
rect 15246 10039 15247 10065
rect 15247 10039 15273 10065
rect 15273 10039 15274 10065
rect 15246 10038 15274 10039
rect 15302 10009 15330 10010
rect 15302 9983 15303 10009
rect 15303 9983 15329 10009
rect 15329 9983 15330 10009
rect 15302 9982 15330 9983
rect 16422 10374 16450 10402
rect 18830 10401 18858 10402
rect 18830 10375 18831 10401
rect 18831 10375 18857 10401
rect 18857 10375 18858 10401
rect 18830 10374 18858 10375
rect 20006 10038 20034 10066
rect 16310 9982 16338 10010
rect 18830 10009 18858 10010
rect 18830 9983 18831 10009
rect 18831 9983 18857 10009
rect 18857 9983 18858 10009
rect 18830 9982 18858 9983
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 9758 20034 9786
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 14966 9086 14994 9114
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14966 8833 14994 8834
rect 14966 8807 14967 8833
rect 14967 8807 14993 8833
rect 14993 8807 14994 8833
rect 14966 8806 14994 8807
rect 15358 8806 15386 8834
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 14686 7910 14714 7938
rect 15022 7910 15050 7938
rect 14798 7601 14826 7602
rect 14798 7575 14799 7601
rect 14799 7575 14825 7601
rect 14825 7575 14826 7601
rect 14798 7574 14826 7575
rect 20006 8414 20034 8442
rect 18830 7574 18858 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 13286 6846 13314 6874
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 12838 2590 12866 2618
rect 12446 2030 12474 2058
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 13398 2617 13426 2618
rect 13398 2591 13399 2617
rect 13399 2591 13425 2617
rect 13425 2591 13426 2617
rect 13398 2590 13426 2591
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 12777 19278 12782 19306
rect 12810 19278 13398 19306
rect 13426 19278 13431 19306
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8409 19110 8414 19138
rect 8442 19110 9030 19138
rect 9058 19110 9063 19138
rect 10425 19110 10430 19138
rect 10458 19110 11046 19138
rect 11074 19110 11079 19138
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 13113 19110 13118 19138
rect 13146 19110 14686 19138
rect 14714 19110 14719 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10089 18718 10094 18746
rect 10122 18718 10710 18746
rect 10738 18718 10743 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 2137 13510 2142 13538
rect 2170 13510 6062 13538
rect 6090 13510 6095 13538
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 12329 13454 12334 13482
rect 12362 13454 13398 13482
rect 13426 13454 13431 13482
rect 0 13440 400 13454
rect 7457 13398 7462 13426
rect 7490 13398 7854 13426
rect 7882 13398 7887 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 12105 13230 12110 13258
rect 12138 13230 12670 13258
rect 12698 13230 12703 13258
rect 13113 13230 13118 13258
rect 13146 13230 14294 13258
rect 14322 13230 14327 13258
rect 7065 13174 7070 13202
rect 7098 13174 7406 13202
rect 7434 13174 7439 13202
rect 8745 13174 8750 13202
rect 8778 13174 10318 13202
rect 10346 13174 10351 13202
rect 10873 13174 10878 13202
rect 10906 13174 12726 13202
rect 12754 13174 12759 13202
rect 0 13146 400 13160
rect 20600 13146 21000 13160
rect 0 13118 966 13146
rect 994 13118 999 13146
rect 10705 13118 10710 13146
rect 10738 13118 11774 13146
rect 11802 13118 12334 13146
rect 12362 13118 12367 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 0 13104 400 13118
rect 20600 13104 21000 13118
rect 6057 13062 6062 13090
rect 6090 13062 7574 13090
rect 7602 13062 7607 13090
rect 14905 13006 14910 13034
rect 14938 13006 15302 13034
rect 15330 13006 18942 13034
rect 18970 13006 18975 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 9305 12838 9310 12866
rect 9338 12838 10710 12866
rect 10738 12838 10743 12866
rect 20600 12810 21000 12824
rect 10145 12782 10150 12810
rect 10178 12782 10822 12810
rect 10850 12782 10855 12810
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 20600 12768 21000 12782
rect 9697 12726 9702 12754
rect 9730 12726 10206 12754
rect 10234 12726 10239 12754
rect 11825 12726 11830 12754
rect 11858 12726 12334 12754
rect 12362 12726 14238 12754
rect 14266 12726 14271 12754
rect 6953 12670 6958 12698
rect 6986 12670 7518 12698
rect 7546 12670 7551 12698
rect 7625 12670 7630 12698
rect 7658 12670 9198 12698
rect 9226 12670 9231 12698
rect 9809 12670 9814 12698
rect 9842 12670 9870 12698
rect 9898 12670 9903 12698
rect 9977 12670 9982 12698
rect 10010 12670 10654 12698
rect 10682 12670 10687 12698
rect 11545 12670 11550 12698
rect 11578 12670 12110 12698
rect 12138 12670 12143 12698
rect 12385 12670 12390 12698
rect 12418 12670 12950 12698
rect 12978 12670 12983 12698
rect 13785 12670 13790 12698
rect 13818 12670 14518 12698
rect 14546 12670 14551 12698
rect 14625 12670 14630 12698
rect 14658 12670 14854 12698
rect 14882 12670 18830 12698
rect 18858 12670 18863 12698
rect 7401 12614 7406 12642
rect 7434 12614 8078 12642
rect 8106 12614 8750 12642
rect 8778 12614 8783 12642
rect 9753 12614 9758 12642
rect 9786 12614 10094 12642
rect 10122 12614 10127 12642
rect 10761 12614 10766 12642
rect 10794 12614 11102 12642
rect 11130 12614 11135 12642
rect 11769 12614 11774 12642
rect 11802 12614 12278 12642
rect 12306 12614 13734 12642
rect 13762 12614 13767 12642
rect 7681 12558 7686 12586
rect 7714 12558 8302 12586
rect 8330 12558 8638 12586
rect 8666 12558 8671 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 8465 12502 8470 12530
rect 8498 12502 9030 12530
rect 9058 12502 9534 12530
rect 9562 12502 9567 12530
rect 0 12474 400 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 6673 12446 6678 12474
rect 6706 12446 7350 12474
rect 7378 12446 7383 12474
rect 7849 12446 7854 12474
rect 7882 12446 7887 12474
rect 9137 12446 9142 12474
rect 9170 12446 10206 12474
rect 10234 12446 10239 12474
rect 0 12432 400 12446
rect 7854 12362 7882 12446
rect 9249 12390 9254 12418
rect 9282 12390 9814 12418
rect 9842 12390 9847 12418
rect 7289 12334 7294 12362
rect 7322 12334 7882 12362
rect 8017 12334 8022 12362
rect 8050 12334 8862 12362
rect 8890 12334 8895 12362
rect 2137 12278 2142 12306
rect 2170 12278 5614 12306
rect 5642 12278 5647 12306
rect 10486 12278 12782 12306
rect 12810 12278 12815 12306
rect 10486 12250 10514 12278
rect 9795 12222 9814 12250
rect 9842 12222 10486 12250
rect 10514 12222 10519 12250
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 10425 12054 10430 12082
rect 10458 12054 11494 12082
rect 11522 12054 11527 12082
rect 5609 11998 5614 12026
rect 5642 11998 7126 12026
rect 7154 11998 7159 12026
rect 13841 11998 13846 12026
rect 13874 11998 14014 12026
rect 14042 11998 14294 12026
rect 14322 11998 14574 12026
rect 14602 11998 15078 12026
rect 15106 11998 15111 12026
rect 15185 11998 15190 12026
rect 15218 11998 16030 12026
rect 16058 11998 18830 12026
rect 18858 11998 18863 12026
rect 8801 11942 8806 11970
rect 8834 11942 9254 11970
rect 9282 11942 9287 11970
rect 11153 11942 11158 11970
rect 11186 11942 11191 11970
rect 11158 11914 11186 11942
rect 9081 11886 9086 11914
rect 9114 11886 9534 11914
rect 9562 11886 9870 11914
rect 9898 11886 9903 11914
rect 10761 11886 10766 11914
rect 10794 11886 11186 11914
rect 8521 11830 8526 11858
rect 8554 11830 9590 11858
rect 9618 11830 9814 11858
rect 9842 11830 9847 11858
rect 9977 11830 9982 11858
rect 10010 11830 10822 11858
rect 10850 11830 11158 11858
rect 11186 11830 11191 11858
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 8913 11718 8918 11746
rect 8946 11718 9842 11746
rect 10089 11718 10094 11746
rect 10122 11718 10654 11746
rect 10682 11718 11326 11746
rect 11354 11718 11359 11746
rect 9814 11690 9842 11718
rect 7681 11662 7686 11690
rect 7714 11662 7910 11690
rect 7938 11662 8862 11690
rect 8890 11662 8895 11690
rect 9814 11662 14798 11690
rect 14826 11662 14831 11690
rect 8969 11606 8974 11634
rect 9002 11606 9534 11634
rect 9562 11606 11410 11634
rect 11489 11606 11494 11634
rect 11522 11606 11830 11634
rect 11858 11606 11863 11634
rect 11382 11578 11410 11606
rect 2137 11550 2142 11578
rect 2170 11550 4214 11578
rect 10537 11550 10542 11578
rect 10570 11550 10990 11578
rect 11018 11550 11023 11578
rect 11382 11550 12054 11578
rect 12082 11550 12087 11578
rect 14681 11550 14686 11578
rect 14714 11550 15246 11578
rect 15274 11550 15279 11578
rect 4186 11522 4214 11550
rect 4186 11494 5614 11522
rect 5642 11494 5647 11522
rect 6673 11494 6678 11522
rect 6706 11494 7406 11522
rect 7434 11494 7439 11522
rect 9753 11494 9758 11522
rect 9786 11494 10262 11522
rect 10290 11494 10710 11522
rect 10738 11494 10743 11522
rect 0 11466 400 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 0 11424 400 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 7625 11270 7630 11298
rect 7658 11270 10598 11298
rect 10626 11270 10631 11298
rect 7849 11214 7854 11242
rect 7882 11214 8022 11242
rect 8050 11214 8055 11242
rect 9025 11214 9030 11242
rect 9058 11214 9534 11242
rect 9562 11214 11998 11242
rect 12026 11214 12031 11242
rect 13337 11214 13342 11242
rect 13370 11214 13790 11242
rect 13818 11214 15974 11242
rect 15946 11186 15974 11214
rect 7233 11158 7238 11186
rect 7266 11158 7798 11186
rect 7826 11158 7831 11186
rect 7961 11158 7966 11186
rect 7994 11158 9702 11186
rect 9730 11158 9735 11186
rect 10369 11158 10374 11186
rect 10402 11158 10542 11186
rect 10570 11158 10575 11186
rect 15946 11158 18830 11186
rect 18858 11158 18863 11186
rect 9702 11130 9730 11158
rect 20600 11130 21000 11144
rect 5609 11102 5614 11130
rect 5642 11102 7182 11130
rect 7210 11102 7215 11130
rect 9702 11102 10822 11130
rect 10850 11102 10855 11130
rect 10985 11102 10990 11130
rect 11018 11102 11494 11130
rect 11522 11102 11527 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 6057 11046 6062 11074
rect 6090 11046 7686 11074
rect 7714 11046 7719 11074
rect 9529 11046 9534 11074
rect 9562 11046 9982 11074
rect 10010 11046 10015 11074
rect 12161 11046 12166 11074
rect 12194 11046 12670 11074
rect 12698 11046 13118 11074
rect 13146 11046 13151 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 8353 10878 8358 10906
rect 8386 10878 9310 10906
rect 9338 10878 9646 10906
rect 9674 10878 9679 10906
rect 11265 10878 11270 10906
rect 11298 10878 11942 10906
rect 11970 10878 11975 10906
rect 13426 10878 14014 10906
rect 14042 10878 14630 10906
rect 14658 10878 14910 10906
rect 14938 10878 14943 10906
rect 13426 10850 13454 10878
rect 7345 10822 7350 10850
rect 7378 10822 8750 10850
rect 8778 10822 9254 10850
rect 9282 10822 9287 10850
rect 10593 10822 10598 10850
rect 10626 10822 10766 10850
rect 10794 10822 10799 10850
rect 12385 10822 12390 10850
rect 12418 10822 12894 10850
rect 12922 10822 13454 10850
rect 20600 10794 21000 10808
rect 11657 10766 11662 10794
rect 11690 10766 12110 10794
rect 12138 10766 12614 10794
rect 12642 10766 12647 10794
rect 15946 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 15946 10738 15974 10766
rect 20600 10752 21000 10766
rect 7121 10710 7126 10738
rect 7154 10710 7462 10738
rect 7490 10710 7495 10738
rect 14065 10710 14070 10738
rect 14098 10710 14350 10738
rect 14378 10710 15974 10738
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 8129 10542 8134 10570
rect 8162 10542 9254 10570
rect 9282 10542 9814 10570
rect 9842 10542 10150 10570
rect 10178 10542 10183 10570
rect 7513 10486 7518 10514
rect 7546 10486 7742 10514
rect 7770 10486 11214 10514
rect 11242 10486 11550 10514
rect 11578 10486 11583 10514
rect 20600 10458 21000 10472
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 20600 10416 21000 10430
rect 8521 10374 8526 10402
rect 8554 10374 9086 10402
rect 9114 10374 9119 10402
rect 11321 10374 11326 10402
rect 11354 10374 11662 10402
rect 11690 10374 11695 10402
rect 16417 10374 16422 10402
rect 16450 10374 18830 10402
rect 18858 10374 18863 10402
rect 10705 10318 10710 10346
rect 10738 10318 10878 10346
rect 10906 10318 10911 10346
rect 9865 10262 9870 10290
rect 9898 10262 11102 10290
rect 11130 10262 11135 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 20600 10122 21000 10136
rect 5665 10094 5670 10122
rect 5698 10094 7238 10122
rect 7266 10094 7271 10122
rect 7681 10094 7686 10122
rect 7714 10094 8078 10122
rect 8106 10094 8111 10122
rect 9179 10094 9198 10122
rect 9226 10094 9231 10122
rect 20006 10094 21000 10122
rect 20006 10066 20034 10094
rect 20600 10080 21000 10094
rect 7345 10038 7350 10066
rect 7378 10038 8134 10066
rect 8162 10038 8167 10066
rect 8241 10038 8246 10066
rect 8274 10038 9758 10066
rect 9786 10038 9791 10066
rect 10817 10038 10822 10066
rect 10850 10038 11494 10066
rect 11522 10038 11527 10066
rect 12670 10038 13398 10066
rect 13426 10038 14126 10066
rect 14154 10038 14406 10066
rect 14434 10038 14439 10066
rect 15241 10038 15246 10066
rect 15274 10038 15974 10066
rect 20001 10038 20006 10066
rect 20034 10038 20039 10066
rect 12670 10010 12698 10038
rect 15946 10010 15974 10038
rect 7625 9982 7630 10010
rect 7658 9982 8302 10010
rect 8330 9982 8335 10010
rect 8633 9982 8638 10010
rect 8666 9982 8918 10010
rect 8946 9982 8951 10010
rect 9361 9982 9366 10010
rect 9394 9982 10374 10010
rect 10402 9982 10407 10010
rect 11153 9982 11158 10010
rect 11186 9982 12698 10010
rect 12777 9982 12782 10010
rect 12810 9982 13230 10010
rect 13258 9982 13678 10010
rect 13706 9982 13711 10010
rect 13897 9982 13902 10010
rect 13930 9982 14238 10010
rect 14266 9982 14271 10010
rect 14681 9982 14686 10010
rect 14714 9982 15302 10010
rect 15330 9982 15335 10010
rect 15946 9982 16310 10010
rect 16338 9982 18830 10010
rect 18858 9982 18863 10010
rect 8969 9926 8974 9954
rect 9002 9926 9310 9954
rect 9338 9926 9343 9954
rect 9417 9926 9422 9954
rect 9450 9926 10598 9954
rect 10626 9926 10631 9954
rect 13449 9926 13454 9954
rect 13482 9926 13958 9954
rect 13986 9926 13991 9954
rect 7737 9870 7742 9898
rect 7770 9870 8806 9898
rect 8834 9870 11550 9898
rect 11578 9870 11583 9898
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 8857 9702 8862 9730
rect 8890 9702 13566 9730
rect 13594 9702 13599 9730
rect 7905 9646 7910 9674
rect 7938 9646 11914 9674
rect 13225 9646 13230 9674
rect 13258 9646 13622 9674
rect 13650 9646 13655 9674
rect 14289 9646 14294 9674
rect 14322 9646 15974 9674
rect 11886 9618 11914 9646
rect 15946 9618 15974 9646
rect 8857 9590 8862 9618
rect 8890 9590 9142 9618
rect 9170 9590 9175 9618
rect 9753 9590 9758 9618
rect 9786 9590 9954 9618
rect 10201 9590 10206 9618
rect 10234 9590 10878 9618
rect 10906 9590 10911 9618
rect 11881 9590 11886 9618
rect 11914 9590 12166 9618
rect 12194 9590 12199 9618
rect 15946 9590 18830 9618
rect 18858 9590 18863 9618
rect 9926 9562 9954 9590
rect 7905 9534 7910 9562
rect 7938 9534 8806 9562
rect 8834 9534 9842 9562
rect 9921 9534 9926 9562
rect 9954 9534 10150 9562
rect 10178 9534 10183 9562
rect 11209 9534 11214 9562
rect 11242 9534 12110 9562
rect 12138 9534 12143 9562
rect 9814 9506 9842 9534
rect 2081 9478 2086 9506
rect 2114 9478 9590 9506
rect 9618 9478 9623 9506
rect 9814 9478 10038 9506
rect 10066 9478 10934 9506
rect 10962 9478 10967 9506
rect 11657 9478 11662 9506
rect 11690 9478 11998 9506
rect 12026 9478 12031 9506
rect 9025 9422 9030 9450
rect 9058 9422 9198 9450
rect 9226 9422 9231 9450
rect 11545 9422 11550 9450
rect 11578 9422 11774 9450
rect 11802 9422 11807 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 7233 9310 7238 9338
rect 7266 9310 7406 9338
rect 7434 9310 7742 9338
rect 7770 9310 7775 9338
rect 10593 9310 10598 9338
rect 10626 9310 12838 9338
rect 12866 9310 12871 9338
rect 5945 9254 5950 9282
rect 5978 9254 8078 9282
rect 8106 9254 8862 9282
rect 8890 9254 8895 9282
rect 11825 9254 11830 9282
rect 11858 9254 12166 9282
rect 12194 9254 12558 9282
rect 12586 9254 12950 9282
rect 12978 9254 12983 9282
rect 9753 9198 9758 9226
rect 9786 9198 9870 9226
rect 9898 9198 10990 9226
rect 11018 9198 11023 9226
rect 12217 9198 12222 9226
rect 12250 9198 12614 9226
rect 12642 9198 12647 9226
rect 13057 9198 13062 9226
rect 13090 9198 14910 9226
rect 14938 9198 14943 9226
rect 7009 9142 7014 9170
rect 7042 9142 7350 9170
rect 7378 9142 7383 9170
rect 8241 9142 8246 9170
rect 8274 9142 9590 9170
rect 9618 9142 9623 9170
rect 9697 9142 9702 9170
rect 9730 9142 10206 9170
rect 10234 9142 10654 9170
rect 10682 9142 10687 9170
rect 13113 9142 13118 9170
rect 13146 9142 13454 9170
rect 13482 9142 13487 9170
rect 9417 9086 9422 9114
rect 9450 9086 11494 9114
rect 11522 9086 11527 9114
rect 13393 9086 13398 9114
rect 13426 9086 14966 9114
rect 14994 9086 14999 9114
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 12497 8974 12502 9002
rect 12530 8974 12782 9002
rect 12810 8974 12815 9002
rect 12665 8918 12670 8946
rect 12698 8918 12703 8946
rect 12670 8890 12698 8918
rect 11321 8862 11326 8890
rect 11354 8862 12334 8890
rect 12362 8862 12698 8890
rect 8801 8806 8806 8834
rect 8834 8806 10710 8834
rect 10738 8806 10743 8834
rect 11489 8806 11494 8834
rect 11522 8806 12950 8834
rect 12978 8806 13398 8834
rect 13426 8806 13431 8834
rect 14961 8806 14966 8834
rect 14994 8806 15358 8834
rect 15386 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 6001 8750 6006 8778
rect 6034 8750 6902 8778
rect 6930 8750 9478 8778
rect 9506 8750 9511 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 9921 8470 9926 8498
rect 9954 8470 11046 8498
rect 11074 8470 11079 8498
rect 13953 8470 13958 8498
rect 13986 8470 14294 8498
rect 14322 8470 14327 8498
rect 20600 8442 21000 8456
rect 8969 8414 8974 8442
rect 9002 8414 9814 8442
rect 9842 8414 9847 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 20600 8400 21000 8414
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 12441 8134 12446 8162
rect 12474 8134 14574 8162
rect 14602 8134 14607 8162
rect 8297 7910 8302 7938
rect 8330 7910 8414 7938
rect 8442 7910 8447 7938
rect 8689 7910 8694 7938
rect 8722 7910 9254 7938
rect 9282 7910 9287 7938
rect 12273 7910 12278 7938
rect 12306 7910 12782 7938
rect 12810 7910 12815 7938
rect 13281 7910 13286 7938
rect 13314 7910 13734 7938
rect 13762 7910 14686 7938
rect 14714 7910 15022 7938
rect 15050 7910 15055 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 8297 7630 8302 7658
rect 8330 7630 8638 7658
rect 8666 7630 8671 7658
rect 7177 7574 7182 7602
rect 7210 7574 8750 7602
rect 8778 7574 8783 7602
rect 12777 7574 12782 7602
rect 12810 7574 13062 7602
rect 13090 7574 13095 7602
rect 14793 7574 14798 7602
rect 14826 7574 18830 7602
rect 18858 7574 18863 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 7233 7350 7238 7378
rect 7266 7350 8470 7378
rect 8498 7350 8503 7378
rect 8577 7350 8582 7378
rect 8610 7350 8974 7378
rect 9002 7350 9310 7378
rect 9338 7350 10878 7378
rect 10906 7350 10911 7378
rect 8241 7294 8246 7322
rect 8274 7294 8694 7322
rect 8722 7294 9086 7322
rect 9114 7294 9119 7322
rect 6897 7238 6902 7266
rect 6930 7238 8358 7266
rect 8386 7238 8806 7266
rect 8834 7238 9310 7266
rect 9338 7238 9343 7266
rect 10201 7238 10206 7266
rect 10234 7238 11270 7266
rect 11298 7238 11303 7266
rect 8969 7182 8974 7210
rect 9002 7182 9254 7210
rect 9282 7182 9287 7210
rect 9641 7126 9646 7154
rect 9674 7126 10710 7154
rect 10738 7126 10743 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 9305 6846 9310 6874
rect 9338 6846 10318 6874
rect 10346 6846 10766 6874
rect 10794 6846 10799 6874
rect 10929 6846 10934 6874
rect 10962 6846 11606 6874
rect 11634 6846 12670 6874
rect 12698 6846 13286 6874
rect 13314 6846 13319 6874
rect 11433 6790 11438 6818
rect 11466 6790 12278 6818
rect 12306 6790 12311 6818
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9809 5054 9814 5082
rect 9842 5054 10206 5082
rect 10234 5054 10239 5082
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 12833 2590 12838 2618
rect 12866 2590 13398 2618
rect 13426 2590 13431 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8073 2086 8078 2114
rect 8106 2086 9254 2114
rect 9282 2086 9287 2114
rect 10089 2030 10094 2058
rect 10122 2030 10710 2058
rect 10738 2030 10743 2058
rect 12441 2030 12446 2058
rect 12474 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10761 1806 10766 1834
rect 10794 1806 11214 1834
rect 11242 1806 11247 1834
rect 11769 1806 11774 1834
rect 11802 1806 12782 1834
rect 12810 1806 12815 1834
rect 8409 1694 8414 1722
rect 8442 1694 9030 1722
rect 9058 1694 9063 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9814 12670 9842 12698
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 9814 12222 9842 12250
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 9198 10094 9226 10122
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9198 9422 9226 9450
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9814 12698 9842 12703
rect 9814 12250 9842 12670
rect 9814 12217 9842 12222
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 9198 10122 9226 10127
rect 9198 9450 9226 10094
rect 9198 9417 9226 9422
rect 9904 9422 10064 10178
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14728 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11312 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 7336 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7448 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11984 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7616 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _123_
timestamp 1698175906
transform 1 0 9632 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _124_
timestamp 1698175906
transform 1 0 10920 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11312 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 7112 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _127_
timestamp 1698175906
transform 1 0 9128 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform 1 0 9296 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12152 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11424 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _132_
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform -1 0 12264 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform -1 0 11760 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _135_
timestamp 1698175906
transform 1 0 12712 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _136_
timestamp 1698175906
transform 1 0 13328 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform 1 0 8008 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9856 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _139_
timestamp 1698175906
transform -1 0 8848 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_
timestamp 1698175906
transform -1 0 9352 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9352 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _142_
timestamp 1698175906
transform -1 0 9968 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 12208 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 11480 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_
timestamp 1698175906
transform -1 0 11088 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9968 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7784 0 -1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _150_
timestamp 1698175906
transform -1 0 7168 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9128 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform 1 0 9632 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform 1 0 10192 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform 1 0 11424 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform 1 0 8120 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform 1 0 9744 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform 1 0 10920 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _159_
timestamp 1698175906
transform -1 0 11480 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _160_
timestamp 1698175906
transform -1 0 11424 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _161_
timestamp 1698175906
transform 1 0 9688 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _162_
timestamp 1698175906
transform 1 0 11256 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _163_
timestamp 1698175906
transform 1 0 11032 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _164_
timestamp 1698175906
transform 1 0 14448 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 15064 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 14392 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _167_
timestamp 1698175906
transform -1 0 8232 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_
timestamp 1698175906
transform 1 0 8176 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _169_
timestamp 1698175906
transform 1 0 8736 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _171_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9128 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform 1 0 9240 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 14784 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform -1 0 13888 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _175_
timestamp 1698175906
transform -1 0 8624 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _176_
timestamp 1698175906
transform -1 0 8064 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9744 0 1 11760
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _178_
timestamp 1698175906
transform 1 0 8008 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _179_
timestamp 1698175906
transform -1 0 8008 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11032 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _181_
timestamp 1698175906
transform -1 0 9912 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _182_
timestamp 1698175906
transform -1 0 10360 0 1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform 1 0 11928 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform -1 0 13496 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _186_
timestamp 1698175906
transform 1 0 12600 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _187_
timestamp 1698175906
transform 1 0 10640 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _188_
timestamp 1698175906
transform -1 0 10864 0 -1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _189_
timestamp 1698175906
transform 1 0 9464 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_
timestamp 1698175906
transform -1 0 15064 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _193_
timestamp 1698175906
transform 1 0 13216 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _194_
timestamp 1698175906
transform 1 0 13720 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _195_
timestamp 1698175906
transform 1 0 11536 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698175906
transform -1 0 11928 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698175906
transform 1 0 12096 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _198_
timestamp 1698175906
transform -1 0 12096 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _199_
timestamp 1698175906
transform 1 0 8736 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _200_
timestamp 1698175906
transform 1 0 8848 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _201_
timestamp 1698175906
transform 1 0 9688 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _202_
timestamp 1698175906
transform -1 0 10024 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _203_
timestamp 1698175906
transform -1 0 9632 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _204_
timestamp 1698175906
transform 1 0 10136 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _205_
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _206_
timestamp 1698175906
transform 1 0 8456 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8120 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _208_
timestamp 1698175906
transform 1 0 8344 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _209_
timestamp 1698175906
transform 1 0 11200 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _210_
timestamp 1698175906
transform -1 0 11704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _211_
timestamp 1698175906
transform 1 0 12712 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _212_
timestamp 1698175906
transform 1 0 12152 0 1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _213_
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _214_
timestamp 1698175906
transform -1 0 14504 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _215_
timestamp 1698175906
transform 1 0 13496 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _216_
timestamp 1698175906
transform 1 0 7056 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _217_
timestamp 1698175906
transform 1 0 7224 0 -1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _218_
timestamp 1698175906
transform -1 0 15400 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _219_
timestamp 1698175906
transform -1 0 15120 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _220_
timestamp 1698175906
transform -1 0 9072 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _221_
timestamp 1698175906
transform -1 0 15344 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _222_
timestamp 1698175906
transform -1 0 14952 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _223_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _224_
timestamp 1698175906
transform 1 0 6888 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _225_
timestamp 1698175906
transform -1 0 7336 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _226_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11256 0 1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _227_
timestamp 1698175906
transform 1 0 7280 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _228_
timestamp 1698175906
transform -1 0 14224 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _229_
timestamp 1698175906
transform 1 0 13048 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13272 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 6720 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 10584 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 13776 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 5488 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 5544 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 8736 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 13328 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 7000 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 8848 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 12264 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 8680 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 13832 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 11536 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 8512 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 9184 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 6776 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _248_
timestamp 1698175906
transform 1 0 10808 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _249_
timestamp 1698175906
transform 1 0 11648 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _250_
timestamp 1698175906
transform 1 0 12768 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _251_
timestamp 1698175906
transform -1 0 7168 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _252_
timestamp 1698175906
transform 1 0 14560 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _253_
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _254_
timestamp 1698175906
transform -1 0 7616 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _255_
timestamp 1698175906
transform -1 0 7168 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _256_
timestamp 1698175906
transform 1 0 12824 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _257_
timestamp 1698175906
transform 1 0 12880 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _258_
timestamp 1698175906
transform 1 0 12712 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _259_
timestamp 1698175906
transform 1 0 16184 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 8344 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 13664 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 7112 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 7280 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 7336 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 10696 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 15064 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 8736 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 10696 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 14000 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 10416 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 13720 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 13272 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform -1 0 10360 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 10808 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 8792 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__CLK
timestamp 1698175906
transform 1 0 13384 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__CLK
timestamp 1698175906
transform 1 0 14616 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__CLK
timestamp 1698175906
transform 1 0 7224 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__CLK
timestamp 1698175906
transform 1 0 14616 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__CLK
timestamp 1698175906
transform 1 0 14280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__CLK
timestamp 1698175906
transform 1 0 8064 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__CLK
timestamp 1698175906
transform 1 0 7392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__CLK
timestamp 1698175906
transform 1 0 14896 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 9632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 11424 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11592 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 10136 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_168
timestamp 1698175906
transform 1 0 10080 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11592 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 12040 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_209
timestamp 1698175906
transform 1 0 12376 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698175906
transform 1 0 14280 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_139
timestamp 1698175906
transform 1 0 8456 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_169
timestamp 1698175906
transform 1 0 10136 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 10360 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_183
timestamp 1698175906
transform 1 0 10920 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_215 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12712 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698175906
transform 1 0 13608 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698175906
transform 1 0 14056 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698175906
transform 1 0 14280 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698175906
transform 1 0 8456 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698175906
transform 1 0 9072 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698175906
transform 1 0 12768 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_143
timestamp 1698175906
transform 1 0 8680 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_147
timestamp 1698175906
transform 1 0 8904 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_151
timestamp 1698175906
transform 1 0 9128 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_160
timestamp 1698175906
transform 1 0 9632 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_167
timestamp 1698175906
transform 1 0 10024 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_187
timestamp 1698175906
transform 1 0 11144 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_223
timestamp 1698175906
transform 1 0 13160 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_227
timestamp 1698175906
transform 1 0 13384 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 14280 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_108
timestamp 1698175906
transform 1 0 6720 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_155
timestamp 1698175906
transform 1 0 9352 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_171
timestamp 1698175906
transform 1 0 10248 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_179
timestamp 1698175906
transform 1 0 10696 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_186
timestamp 1698175906
transform 1 0 11088 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_188
timestamp 1698175906
transform 1 0 11200 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_197
timestamp 1698175906
transform 1 0 11704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698175906
transform 1 0 12152 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_221
timestamp 1698175906
transform 1 0 13048 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_254
timestamp 1698175906
transform 1 0 14896 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_258
timestamp 1698175906
transform 1 0 15120 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698175906
transform 1 0 16016 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 16240 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_123
timestamp 1698175906
transform 1 0 7560 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_131
timestamp 1698175906
transform 1 0 8008 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_156
timestamp 1698175906
transform 1 0 9408 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_193
timestamp 1698175906
transform 1 0 11480 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_195
timestamp 1698175906
transform 1 0 11592 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_210
timestamp 1698175906
transform 1 0 12432 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_226
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_230
timestamp 1698175906
transform 1 0 13552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_232
timestamp 1698175906
transform 1 0 13664 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_235
timestamp 1698175906
transform 1 0 13832 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 14280 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_251
timestamp 1698175906
transform 1 0 14728 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 5152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698175906
transform 1 0 5376 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_86
timestamp 1698175906
transform 1 0 5488 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_116
timestamp 1698175906
transform 1 0 7168 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_120
timestamp 1698175906
transform 1 0 7392 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 8288 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_158
timestamp 1698175906
transform 1 0 9520 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_160
timestamp 1698175906
transform 1 0 9632 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_167
timestamp 1698175906
transform 1 0 10024 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_199
timestamp 1698175906
transform 1 0 11816 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698175906
transform 1 0 12992 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_224
timestamp 1698175906
transform 1 0 13216 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_232
timestamp 1698175906
transform 1 0 13664 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_234
timestamp 1698175906
transform 1 0 13776 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_264
timestamp 1698175906
transform 1 0 15456 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_109
timestamp 1698175906
transform 1 0 6776 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_116
timestamp 1698175906
transform 1 0 7168 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_132
timestamp 1698175906
transform 1 0 8064 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_140
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 10360 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_181
timestamp 1698175906
transform 1 0 10808 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698175906
transform 1 0 11032 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_187
timestamp 1698175906
transform 1 0 11144 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_193
timestamp 1698175906
transform 1 0 11480 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_199
timestamp 1698175906
transform 1 0 11816 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_203
timestamp 1698175906
transform 1 0 12040 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_225
timestamp 1698175906
transform 1 0 13272 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_239
timestamp 1698175906
transform 1 0 14056 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 14280 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_251
timestamp 1698175906
transform 1 0 14728 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_257
timestamp 1698175906
transform 1 0 15064 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_289
timestamp 1698175906
transform 1 0 16856 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_305
timestamp 1698175906
transform 1 0 17752 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698175906
transform 1 0 18200 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698175906
transform 1 0 5376 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_127
timestamp 1698175906
transform 1 0 7784 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 8232 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_152
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_176
timestamp 1698175906
transform 1 0 10528 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_191
timestamp 1698175906
transform 1 0 11368 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_198
timestamp 1698175906
transform 1 0 11760 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_234
timestamp 1698175906
transform 1 0 13776 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_266
timestamp 1698175906
transform 1 0 15568 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 16016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_117
timestamp 1698175906
transform 1 0 7224 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_135
timestamp 1698175906
transform 1 0 8232 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_143
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_155
timestamp 1698175906
transform 1 0 9352 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_157
timestamp 1698175906
transform 1 0 9464 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698175906
transform 1 0 10304 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_207
timestamp 1698175906
transform 1 0 12264 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_215
timestamp 1698175906
transform 1 0 12712 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_251
timestamp 1698175906
transform 1 0 14728 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_112
timestamp 1698175906
transform 1 0 6944 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_114
timestamp 1698175906
transform 1 0 7056 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 8344 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 8456 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_218
timestamp 1698175906
transform 1 0 12880 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_220
timestamp 1698175906
transform 1 0 12992 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_247
timestamp 1698175906
transform 1 0 14504 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_251
timestamp 1698175906
transform 1 0 14728 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_263
timestamp 1698175906
transform 1 0 15400 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 16296 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698175906
transform 1 0 7112 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_119
timestamp 1698175906
transform 1 0 7336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_132
timestamp 1698175906
transform 1 0 8064 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_147
timestamp 1698175906
transform 1 0 8904 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_159
timestamp 1698175906
transform 1 0 9576 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_283
timestamp 1698175906
transform 1 0 16520 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_117
timestamp 1698175906
transform 1 0 7224 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_121
timestamp 1698175906
transform 1 0 7448 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_129
timestamp 1698175906
transform 1 0 7896 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_133
timestamp 1698175906
transform 1 0 8120 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_197
timestamp 1698175906
transform 1 0 11704 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_199
timestamp 1698175906
transform 1 0 11816 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 12208 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_216
timestamp 1698175906
transform 1 0 12768 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_252
timestamp 1698175906
transform 1 0 14784 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_256
timestamp 1698175906
transform 1 0 15008 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_272
timestamp 1698175906
transform 1 0 15904 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 6888 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_113
timestamp 1698175906
transform 1 0 7000 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_119
timestamp 1698175906
transform 1 0 7336 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_133
timestamp 1698175906
transform 1 0 8120 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_141
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_195
timestamp 1698175906
transform 1 0 11592 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_199
timestamp 1698175906
transform 1 0 11816 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_206
timestamp 1698175906
transform 1 0 12208 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_236
timestamp 1698175906
transform 1 0 13888 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_240
timestamp 1698175906
transform 1 0 14112 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 5152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_84
timestamp 1698175906
transform 1 0 5376 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_86
timestamp 1698175906
transform 1 0 5488 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_116
timestamp 1698175906
transform 1 0 7168 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_132
timestamp 1698175906
transform 1 0 8064 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_152
timestamp 1698175906
transform 1 0 9184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_166
timestamp 1698175906
transform 1 0 9968 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_182
timestamp 1698175906
transform 1 0 10864 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_189
timestamp 1698175906
transform 1 0 11256 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_193
timestamp 1698175906
transform 1 0 11480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_195
timestamp 1698175906
transform 1 0 11592 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_201
timestamp 1698175906
transform 1 0 11928 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_221
timestamp 1698175906
transform 1 0 13048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_223
timestamp 1698175906
transform 1 0 13160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_229
timestamp 1698175906
transform 1 0 13496 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_245
timestamp 1698175906
transform 1 0 14392 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_249
timestamp 1698175906
transform 1 0 14616 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_255
timestamp 1698175906
transform 1 0 14952 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_262
timestamp 1698175906
transform 1 0 15344 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 16240 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698175906
transform 1 0 6888 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_113
timestamp 1698175906
transform 1 0 7000 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_118
timestamp 1698175906
transform 1 0 7280 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_122
timestamp 1698175906
transform 1 0 7504 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_130
timestamp 1698175906
transform 1 0 7952 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_134
timestamp 1698175906
transform 1 0 8176 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_142
timestamp 1698175906
transform 1 0 8624 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_146
timestamp 1698175906
transform 1 0 8848 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_167
timestamp 1698175906
transform 1 0 10024 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_193
timestamp 1698175906
transform 1 0 11480 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_225
timestamp 1698175906
transform 1 0 13272 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_276
timestamp 1698175906
transform 1 0 16128 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_308
timestamp 1698175906
transform 1 0 17920 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698175906
transform 1 0 18144 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698175906
transform 1 0 18256 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 5152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 5376 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698175906
transform 1 0 5488 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_116
timestamp 1698175906
transform 1 0 7168 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_127
timestamp 1698175906
transform 1 0 7784 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 8232 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_158
timestamp 1698175906
transform 1 0 9520 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_173
timestamp 1698175906
transform 1 0 10360 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698175906
transform 1 0 12152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_228
timestamp 1698175906
transform 1 0 13440 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_263
timestamp 1698175906
transform 1 0 15400 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_119
timestamp 1698175906
transform 1 0 7336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_130
timestamp 1698175906
transform 1 0 7952 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_134
timestamp 1698175906
transform 1 0 8176 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_150
timestamp 1698175906
transform 1 0 9072 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_154
timestamp 1698175906
transform 1 0 9296 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_156
timestamp 1698175906
transform 1 0 9408 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698175906
transform 1 0 10360 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_183
timestamp 1698175906
transform 1 0 10920 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_197
timestamp 1698175906
transform 1 0 11704 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_220
timestamp 1698175906
transform 1 0 12992 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_228
timestamp 1698175906
transform 1 0 13440 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_230
timestamp 1698175906
transform 1 0 13552 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_236
timestamp 1698175906
transform 1 0 13888 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_257
timestamp 1698175906
transform 1 0 15064 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_289
timestamp 1698175906
transform 1 0 16856 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_305
timestamp 1698175906
transform 1 0 17752 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698175906
transform 1 0 18200 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_92
timestamp 1698175906
transform 1 0 5824 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_94
timestamp 1698175906
transform 1 0 5936 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_124
timestamp 1698175906
transform 1 0 7616 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_172
timestamp 1698175906
transform 1 0 10304 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_176
timestamp 1698175906
transform 1 0 10528 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_206
timestamp 1698175906
transform 1 0 12208 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_224
timestamp 1698175906
transform 1 0 13216 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_255
timestamp 1698175906
transform 1 0 14952 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_259
timestamp 1698175906
transform 1 0 15176 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_275
timestamp 1698175906
transform 1 0 16072 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 2240 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 2464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_142
timestamp 1698175906
transform 1 0 8624 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_181
timestamp 1698175906
transform 1 0 10808 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_189
timestamp 1698175906
transform 1 0 11256 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_193
timestamp 1698175906
transform 1 0 11480 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_195
timestamp 1698175906
transform 1 0 11592 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_225
timestamp 1698175906
transform 1 0 13272 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_229
timestamp 1698175906
transform 1 0 13496 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_158
timestamp 1698175906
transform 1 0 9520 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_166
timestamp 1698175906
transform 1 0 9968 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 10080 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 11592 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 12040 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 14280 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 16072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_165
timestamp 1698175906
transform 1 0 9912 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 10136 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 10416 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 11928 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 12040 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_266
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 2240 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 8456 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 10136 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 12824 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 12824 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 10136 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 10472 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 8456 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 13104 20600 13160 21000 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 12768 0 12824 400 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 8064 0 8120 400 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 8988 6860 8988 6860 0 _000_
rlabel metal2 9660 7028 9660 7028 0 _001_
rlabel metal2 8484 7336 8484 7336 0 _002_
rlabel metal2 11256 6916 11256 6916 0 _003_
rlabel metal3 12404 13244 12404 13244 0 _004_
rlabel metal2 13636 9800 13636 9800 0 _005_
rlabel metal2 6692 12432 6692 12432 0 _006_
rlabel metal2 14868 10220 14868 10220 0 _007_
rlabel metal2 14700 11788 14700 11788 0 _008_
rlabel metal2 7028 12964 7028 12964 0 _009_
rlabel metal3 7056 11508 7056 11508 0 _010_
rlabel metal2 13188 10416 13188 10416 0 _011_
rlabel metal2 13664 7700 13664 7700 0 _012_
rlabel metal2 7196 7448 7196 7448 0 _013_
rlabel metal2 11284 12936 11284 12936 0 _014_
rlabel metal2 14224 12404 14224 12404 0 _015_
rlabel metal2 8092 9380 8092 9380 0 _016_
rlabel metal2 6020 8624 6020 8624 0 _017_
rlabel metal2 6076 10948 6076 10948 0 _018_
rlabel metal2 9212 8988 9212 8988 0 _019_
rlabel metal2 13776 12852 13776 12852 0 _020_
rlabel metal2 7476 13440 7476 13440 0 _021_
rlabel metal2 10724 12824 10724 12824 0 _022_
rlabel metal2 12740 11368 12740 11368 0 _023_
rlabel metal2 10276 12432 10276 12432 0 _024_
rlabel metal3 14140 8484 14140 8484 0 _025_
rlabel metal2 11984 7308 11984 7308 0 _026_
rlabel metal2 10668 11704 10668 11704 0 _027_
rlabel metal2 14252 12712 14252 12712 0 _028_
rlabel metal2 14532 10430 14532 10430 0 _029_
rlabel metal3 14980 11564 14980 11564 0 _030_
rlabel metal2 14308 12768 14308 12768 0 _031_
rlabel metal2 9268 12180 9268 12180 0 _032_
rlabel metal2 7924 11424 7924 11424 0 _033_
rlabel metal2 9324 9604 9324 9604 0 _034_
rlabel metal3 14168 12684 14168 12684 0 _035_
rlabel metal2 7476 12600 7476 12600 0 _036_
rlabel metal2 7868 12936 7868 12936 0 _037_
rlabel metal2 9016 12348 9016 12348 0 _038_
rlabel metal2 8036 13020 8036 13020 0 _039_
rlabel metal2 12796 12180 12796 12180 0 _040_
rlabel metal2 9772 12544 9772 12544 0 _041_
rlabel metal3 10332 12684 10332 12684 0 _042_
rlabel metal3 12656 11060 12656 11060 0 _043_
rlabel metal2 13132 11564 13132 11564 0 _044_
rlabel metal2 10808 12012 10808 12012 0 _045_
rlabel metal2 10668 11340 10668 11340 0 _046_
rlabel metal2 9996 12236 9996 12236 0 _047_
rlabel metal2 14924 9072 14924 9072 0 _048_
rlabel metal2 13468 9184 13468 9184 0 _049_
rlabel metal2 13804 8960 13804 8960 0 _050_
rlabel metal2 11788 8428 11788 8428 0 _051_
rlabel metal2 11816 8036 11816 8036 0 _052_
rlabel metal2 12012 7952 12012 7952 0 _053_
rlabel metal2 13580 9856 13580 9856 0 _054_
rlabel metal2 9436 7462 9436 7462 0 _055_
rlabel metal3 10752 7252 10752 7252 0 _056_
rlabel metal2 9772 7280 9772 7280 0 _057_
rlabel metal2 10388 7280 10388 7280 0 _058_
rlabel metal2 8316 8568 8316 8568 0 _059_
rlabel metal2 8400 7812 8400 7812 0 _060_
rlabel metal2 11508 7364 11508 7364 0 _061_
rlabel metal3 12684 12684 12684 12684 0 _062_
rlabel metal2 12628 12936 12628 12936 0 _063_
rlabel metal3 14084 9996 14084 9996 0 _064_
rlabel metal2 7280 12068 7280 12068 0 _065_
rlabel metal2 15092 9996 15092 9996 0 _066_
rlabel metal3 9828 11704 9828 11704 0 _067_
rlabel metal2 14980 11564 14980 11564 0 _068_
rlabel metal3 7252 12684 7252 12684 0 _069_
rlabel metal2 7196 11312 7196 11312 0 _070_
rlabel metal2 10640 11060 10640 11060 0 _071_
rlabel metal2 13972 9968 13972 9968 0 _072_
rlabel metal2 12460 8428 12460 8428 0 _073_
rlabel metal2 10836 10220 10836 10220 0 _074_
rlabel metal2 7532 11340 7532 11340 0 _075_
rlabel metal2 8316 10836 8316 10836 0 _076_
rlabel metal3 12040 9604 12040 9604 0 _077_
rlabel metal3 12404 9268 12404 9268 0 _078_
rlabel metal3 8372 9548 8372 9548 0 _079_
rlabel metal2 8008 10444 8008 10444 0 _080_
rlabel metal3 10444 9212 10444 9212 0 _081_
rlabel metal2 11116 10332 11116 10332 0 _082_
rlabel metal2 11340 9156 11340 9156 0 _083_
rlabel metal2 10164 10444 10164 10444 0 _084_
rlabel metal2 9380 12152 9380 12152 0 _085_
rlabel metal3 9268 11620 9268 11620 0 _086_
rlabel metal2 12796 8904 12796 8904 0 _087_
rlabel metal2 7756 10808 7756 10808 0 _088_
rlabel metal3 12376 10780 12376 10780 0 _089_
rlabel metal2 13300 9128 13300 9128 0 _090_
rlabel metal2 11676 9352 11676 9352 0 _091_
rlabel metal2 14980 9576 14980 9576 0 _092_
rlabel metal2 13412 8596 13412 8596 0 _093_
rlabel metal2 8260 10248 8260 10248 0 _094_
rlabel metal2 9828 9044 9828 9044 0 _095_
rlabel metal3 8988 7924 8988 7924 0 _096_
rlabel metal2 8876 7728 8876 7728 0 _097_
rlabel metal2 12012 11200 12012 11200 0 _098_
rlabel metal3 8932 9156 8932 9156 0 _099_
rlabel metal3 8428 12684 8428 12684 0 _100_
rlabel metal2 11284 11704 11284 11704 0 _101_
rlabel metal2 11340 7644 11340 7644 0 _102_
rlabel metal3 9156 7364 9156 7364 0 _103_
rlabel metal2 10332 10388 10332 10388 0 _104_
rlabel metal2 7084 8988 7084 8988 0 _105_
rlabel metal2 10780 11004 10780 11004 0 _106_
rlabel metal2 9772 10948 9772 10948 0 _107_
rlabel metal2 10444 11872 10444 11872 0 _108_
rlabel metal2 11480 12852 11480 12852 0 _109_
rlabel metal2 9548 11956 9548 11956 0 _110_
rlabel metal3 10416 11844 10416 11844 0 _111_
rlabel metal2 10556 11396 10556 11396 0 _112_
rlabel metal2 12292 12656 12292 12656 0 _113_
rlabel metal2 11116 12404 11116 12404 0 _114_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 11676 10220 11676 10220 0 clknet_0_clk
rlabel metal2 10332 6692 10332 6692 0 clknet_1_0__leaf_clk
rlabel metal3 12880 13468 12880 13468 0 clknet_1_1__leaf_clk
rlabel metal2 7420 9184 7420 9184 0 dut52.count\[0\]
rlabel metal2 7252 8792 7252 8792 0 dut52.count\[1\]
rlabel metal2 7476 10556 7476 10556 0 dut52.count\[2\]
rlabel metal3 9968 9156 9968 9156 0 dut52.count\[3\]
rlabel metal2 16100 10416 16100 10416 0 net1
rlabel metal2 10696 1764 10696 1764 0 net10
rlabel metal2 12180 15960 12180 15960 0 net11
rlabel metal2 15372 8596 15372 8596 0 net12
rlabel metal2 12908 3374 12908 3374 0 net13
rlabel metal2 12628 4858 12628 4858 0 net14
rlabel metal2 10220 12908 10220 12908 0 net15
rlabel metal2 14364 9856 14364 9856 0 net16
rlabel metal2 2156 12516 2156 12516 0 net17
rlabel metal3 14882 11228 14882 11228 0 net18
rlabel metal2 10332 13580 10332 13580 0 net19
rlabel metal2 6076 13300 6076 13300 0 net2
rlabel metal2 14868 12880 14868 12880 0 net20
rlabel metal2 14924 12852 14924 12852 0 net21
rlabel metal3 8484 7308 8484 7308 0 net22
rlabel metal2 14644 7784 14644 7784 0 net23
rlabel metal2 16436 10360 16436 10360 0 net24
rlabel metal2 8484 13580 8484 13580 0 net25
rlabel metal3 14224 10724 14224 10724 0 net26
rlabel metal2 8316 7616 8316 7616 0 net3
rlabel metal2 12320 6804 12320 6804 0 net4
rlabel metal3 3178 11564 3178 11564 0 net5
rlabel metal2 14308 16128 14308 16128 0 net6
rlabel metal2 10220 3612 10220 3612 0 net7
rlabel metal2 15204 11844 15204 11844 0 net8
rlabel metal2 13104 13580 13104 13580 0 net9
rlabel metal3 20321 10108 20321 10108 0 segm[0]
rlabel metal3 679 13132 679 13132 0 segm[10]
rlabel metal2 8428 1043 8428 1043 0 segm[11]
rlabel metal2 11788 1099 11788 1099 0 segm[12]
rlabel metal3 679 11452 679 11452 0 segm[13]
rlabel metal2 13132 19873 13132 19873 0 segm[1]
rlabel metal2 10108 1211 10108 1211 0 segm[2]
rlabel metal2 20020 12180 20020 12180 0 segm[3]
rlabel metal2 12796 19957 12796 19957 0 segm[4]
rlabel metal2 10780 1099 10780 1099 0 segm[5]
rlabel metal2 12124 19873 12124 19873 0 segm[6]
rlabel metal2 20020 8820 20020 8820 0 segm[7]
rlabel metal2 12796 791 12796 791 0 segm[8]
rlabel metal2 12460 1211 12460 1211 0 segm[9]
rlabel metal2 10108 19677 10108 19677 0 sel[0]
rlabel metal2 20020 9744 20020 9744 0 sel[10]
rlabel metal3 679 12460 679 12460 0 sel[11]
rlabel metal2 20020 11172 20020 11172 0 sel[1]
rlabel metal2 10444 19873 10444 19873 0 sel[2]
rlabel metal2 20020 12908 20020 12908 0 sel[3]
rlabel metal2 20020 13356 20020 13356 0 sel[4]
rlabel metal2 8092 1239 8092 1239 0 sel[5]
rlabel metal2 20020 8400 20020 8400 0 sel[6]
rlabel metal3 20321 10444 20321 10444 0 sel[7]
rlabel metal2 8428 19873 8428 19873 0 sel[8]
rlabel metal2 20020 10752 20020 10752 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
