magic
tech gf180mcuD
magscale 1 10
timestamp 1699641113
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 26126 38274 26178 38286
rect 26126 38210 26178 38222
rect 18834 38110 18846 38162
rect 18898 38110 18910 38162
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 23538 37998 23550 38050
rect 23602 37998 23614 38050
rect 25554 37998 25566 38050
rect 25618 37998 25630 38050
rect 30494 37938 30546 37950
rect 30494 37874 30546 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 22766 37490 22818 37502
rect 22766 37426 22818 37438
rect 26798 37490 26850 37502
rect 26798 37426 26850 37438
rect 20962 37214 20974 37266
rect 21026 37214 21038 37266
rect 22194 37214 22206 37266
rect 22258 37214 22270 37266
rect 25890 37214 25902 37266
rect 25954 37214 25966 37266
rect 19506 37102 19518 37154
rect 19570 37102 19582 37154
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 16718 36706 16770 36718
rect 16718 36642 16770 36654
rect 15698 36430 15710 36482
rect 15762 36430 15774 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 22878 28082 22930 28094
rect 22530 28030 22542 28082
rect 22594 28030 22606 28082
rect 22878 28018 22930 28030
rect 23774 27970 23826 27982
rect 23774 27906 23826 27918
rect 23662 27858 23714 27870
rect 19282 27806 19294 27858
rect 19346 27806 19358 27858
rect 23662 27794 23714 27806
rect 17838 27746 17890 27758
rect 17838 27682 17890 27694
rect 19070 27746 19122 27758
rect 20066 27694 20078 27746
rect 20130 27694 20142 27746
rect 22194 27694 22206 27746
rect 22258 27694 22270 27746
rect 19070 27682 19122 27694
rect 17726 27634 17778 27646
rect 17726 27570 17778 27582
rect 23774 27634 23826 27646
rect 23774 27570 23826 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 1934 27186 1986 27198
rect 16930 27134 16942 27186
rect 16994 27134 17006 27186
rect 19058 27134 19070 27186
rect 19122 27134 19134 27186
rect 23762 27134 23774 27186
rect 23826 27134 23838 27186
rect 25890 27134 25902 27186
rect 25954 27134 25966 27186
rect 1934 27122 1986 27134
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 16146 27022 16158 27074
rect 16210 27022 16222 27074
rect 22978 27022 22990 27074
rect 23042 27022 23054 27074
rect 14254 26962 14306 26974
rect 14254 26898 14306 26910
rect 14366 26962 14418 26974
rect 14366 26898 14418 26910
rect 19518 26962 19570 26974
rect 19518 26898 19570 26910
rect 19630 26962 19682 26974
rect 19630 26898 19682 26910
rect 19294 26850 19346 26862
rect 19294 26786 19346 26798
rect 20078 26850 20130 26862
rect 20078 26786 20130 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 20862 26514 20914 26526
rect 20862 26450 20914 26462
rect 21422 26514 21474 26526
rect 21422 26450 21474 26462
rect 23886 26514 23938 26526
rect 23886 26450 23938 26462
rect 24558 26514 24610 26526
rect 24558 26450 24610 26462
rect 20750 26402 20802 26414
rect 13346 26350 13358 26402
rect 13410 26350 13422 26402
rect 20750 26338 20802 26350
rect 15934 26290 15986 26302
rect 12674 26238 12686 26290
rect 12738 26238 12750 26290
rect 15934 26226 15986 26238
rect 16046 26290 16098 26302
rect 16046 26226 16098 26238
rect 16158 26290 16210 26302
rect 16158 26226 16210 26238
rect 16270 26290 16322 26302
rect 16270 26226 16322 26238
rect 16382 26290 16434 26302
rect 23662 26290 23714 26302
rect 17378 26238 17390 26290
rect 17442 26238 17454 26290
rect 23426 26238 23438 26290
rect 23490 26238 23502 26290
rect 16382 26226 16434 26238
rect 23662 26226 23714 26238
rect 23998 26290 24050 26302
rect 23998 26226 24050 26238
rect 24446 26290 24498 26302
rect 24446 26226 24498 26238
rect 22990 26178 23042 26190
rect 15474 26126 15486 26178
rect 15538 26126 15550 26178
rect 18162 26126 18174 26178
rect 18226 26126 18238 26178
rect 20290 26126 20302 26178
rect 20354 26126 20366 26178
rect 22990 26114 23042 26126
rect 23774 26178 23826 26190
rect 23774 26114 23826 26126
rect 20862 26066 20914 26078
rect 20862 26002 20914 26014
rect 23102 26066 23154 26078
rect 23102 26002 23154 26014
rect 24558 26066 24610 26078
rect 24558 26002 24610 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 19406 25730 19458 25742
rect 15474 25678 15486 25730
rect 15538 25727 15550 25730
rect 15922 25727 15934 25730
rect 15538 25681 15934 25727
rect 15538 25678 15550 25681
rect 15922 25678 15934 25681
rect 15986 25678 15998 25730
rect 19406 25666 19458 25678
rect 22430 25730 22482 25742
rect 22430 25666 22482 25678
rect 13470 25618 13522 25630
rect 14578 25566 14590 25618
rect 14642 25566 14654 25618
rect 16258 25566 16270 25618
rect 16322 25566 16334 25618
rect 20178 25566 20190 25618
rect 20242 25566 20254 25618
rect 23650 25566 23662 25618
rect 23714 25566 23726 25618
rect 25778 25566 25790 25618
rect 25842 25566 25854 25618
rect 13470 25554 13522 25566
rect 14702 25506 14754 25518
rect 17726 25506 17778 25518
rect 17490 25454 17502 25506
rect 17554 25454 17566 25506
rect 14702 25442 14754 25454
rect 17726 25442 17778 25454
rect 17950 25506 18002 25518
rect 17950 25442 18002 25454
rect 18174 25506 18226 25518
rect 18174 25442 18226 25454
rect 18622 25506 18674 25518
rect 18622 25442 18674 25454
rect 18846 25506 18898 25518
rect 18846 25442 18898 25454
rect 19854 25506 19906 25518
rect 20626 25454 20638 25506
rect 20690 25454 20702 25506
rect 22866 25454 22878 25506
rect 22930 25454 22942 25506
rect 19854 25442 19906 25454
rect 15150 25394 15202 25406
rect 15150 25330 15202 25342
rect 16270 25394 16322 25406
rect 16270 25330 16322 25342
rect 16494 25394 16546 25406
rect 16494 25330 16546 25342
rect 17278 25394 17330 25406
rect 17278 25330 17330 25342
rect 19182 25394 19234 25406
rect 19182 25330 19234 25342
rect 20078 25394 20130 25406
rect 20078 25330 20130 25342
rect 20190 25394 20242 25406
rect 20190 25330 20242 25342
rect 22430 25394 22482 25406
rect 22430 25330 22482 25342
rect 22542 25394 22594 25406
rect 22542 25330 22594 25342
rect 13582 25282 13634 25294
rect 13582 25218 13634 25230
rect 14590 25282 14642 25294
rect 14590 25218 14642 25230
rect 14926 25282 14978 25294
rect 14926 25218 14978 25230
rect 15710 25282 15762 25294
rect 15710 25218 15762 25230
rect 17726 25282 17778 25294
rect 17726 25218 17778 25230
rect 18510 25282 18562 25294
rect 18510 25218 18562 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 20402 24894 20414 24946
rect 20466 24894 20478 24946
rect 22642 24894 22654 24946
rect 22706 24894 22718 24946
rect 18398 24834 18450 24846
rect 13906 24782 13918 24834
rect 13970 24782 13982 24834
rect 18398 24770 18450 24782
rect 15150 24722 15202 24734
rect 14578 24670 14590 24722
rect 14642 24670 14654 24722
rect 15150 24658 15202 24670
rect 18734 24722 18786 24734
rect 20750 24722 20802 24734
rect 18946 24670 18958 24722
rect 19010 24670 19022 24722
rect 18734 24658 18786 24670
rect 20750 24658 20802 24670
rect 22318 24722 22370 24734
rect 26562 24670 26574 24722
rect 26626 24670 26638 24722
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 22318 24658 22370 24670
rect 11778 24558 11790 24610
rect 11842 24558 11854 24610
rect 27346 24558 27358 24610
rect 27410 24558 27422 24610
rect 29474 24558 29486 24610
rect 29538 24558 29550 24610
rect 18510 24498 18562 24510
rect 18510 24434 18562 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 27470 24162 27522 24174
rect 27470 24098 27522 24110
rect 40014 24050 40066 24062
rect 40014 23986 40066 23998
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 18510 23826 18562 23838
rect 22654 23826 22706 23838
rect 19282 23774 19294 23826
rect 19346 23774 19358 23826
rect 18510 23762 18562 23774
rect 22654 23762 22706 23774
rect 27582 23826 27634 23838
rect 27582 23762 27634 23774
rect 28030 23826 28082 23838
rect 28030 23762 28082 23774
rect 28254 23826 28306 23838
rect 28254 23762 28306 23774
rect 28366 23826 28418 23838
rect 28366 23762 28418 23774
rect 14366 23714 14418 23726
rect 14366 23650 14418 23662
rect 18622 23714 18674 23726
rect 18622 23650 18674 23662
rect 18958 23714 19010 23726
rect 18958 23650 19010 23662
rect 22542 23714 22594 23726
rect 22542 23650 22594 23662
rect 27470 23714 27522 23726
rect 27470 23650 27522 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 19618 23326 19630 23378
rect 19682 23326 19694 23378
rect 20850 23326 20862 23378
rect 20914 23326 20926 23378
rect 17390 23266 17442 23278
rect 12002 23214 12014 23266
rect 12066 23214 12078 23266
rect 19170 23214 19182 23266
rect 19234 23214 19246 23266
rect 19954 23214 19966 23266
rect 20018 23214 20030 23266
rect 17390 23202 17442 23214
rect 17726 23154 17778 23166
rect 11330 23102 11342 23154
rect 11394 23102 11406 23154
rect 14914 23102 14926 23154
rect 14978 23102 14990 23154
rect 18162 23102 18174 23154
rect 18226 23102 18238 23154
rect 19058 23102 19070 23154
rect 19122 23102 19134 23154
rect 20626 23102 20638 23154
rect 20690 23102 20702 23154
rect 21858 23102 21870 23154
rect 21922 23102 21934 23154
rect 27122 23102 27134 23154
rect 27186 23102 27198 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 17726 23090 17778 23102
rect 14478 23042 14530 23054
rect 18622 23042 18674 23054
rect 14130 22990 14142 23042
rect 14194 22990 14206 23042
rect 15362 22990 15374 23042
rect 15426 22990 15438 23042
rect 22530 22990 22542 23042
rect 22594 22990 22606 23042
rect 24658 22990 24670 23042
rect 24722 22990 24734 23042
rect 27906 22990 27918 23042
rect 27970 22990 27982 23042
rect 30034 22990 30046 23042
rect 30098 22990 30110 23042
rect 14478 22978 14530 22990
rect 18622 22978 18674 22990
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 15150 22594 15202 22606
rect 15150 22530 15202 22542
rect 28478 22594 28530 22606
rect 28478 22530 28530 22542
rect 16382 22482 16434 22494
rect 16382 22418 16434 22430
rect 18958 22482 19010 22494
rect 18958 22418 19010 22430
rect 21310 22482 21362 22494
rect 21310 22418 21362 22430
rect 28590 22482 28642 22494
rect 28590 22418 28642 22430
rect 29262 22482 29314 22494
rect 29262 22418 29314 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 14254 22370 14306 22382
rect 14254 22306 14306 22318
rect 14926 22370 14978 22382
rect 14926 22306 14978 22318
rect 16158 22370 16210 22382
rect 22318 22370 22370 22382
rect 17378 22318 17390 22370
rect 17442 22318 17454 22370
rect 19170 22318 19182 22370
rect 19234 22318 19246 22370
rect 16158 22306 16210 22318
rect 22318 22306 22370 22318
rect 23438 22370 23490 22382
rect 23438 22306 23490 22318
rect 23662 22370 23714 22382
rect 23662 22306 23714 22318
rect 24446 22370 24498 22382
rect 24446 22306 24498 22318
rect 27694 22370 27746 22382
rect 27694 22306 27746 22318
rect 28142 22370 28194 22382
rect 28142 22306 28194 22318
rect 29038 22370 29090 22382
rect 29038 22306 29090 22318
rect 29486 22370 29538 22382
rect 29486 22306 29538 22318
rect 29598 22370 29650 22382
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 29598 22306 29650 22318
rect 17838 22258 17890 22270
rect 17838 22194 17890 22206
rect 20190 22258 20242 22270
rect 22990 22258 23042 22270
rect 23886 22258 23938 22270
rect 21634 22206 21646 22258
rect 21698 22206 21710 22258
rect 22642 22206 22654 22258
rect 22706 22206 22718 22258
rect 23202 22206 23214 22258
rect 23266 22206 23278 22258
rect 20190 22194 20242 22206
rect 22990 22194 23042 22206
rect 23886 22194 23938 22206
rect 24222 22258 24274 22270
rect 24222 22194 24274 22206
rect 24782 22258 24834 22270
rect 24782 22194 24834 22206
rect 27358 22258 27410 22270
rect 27358 22194 27410 22206
rect 27470 22258 27522 22270
rect 27470 22194 27522 22206
rect 13918 22146 13970 22158
rect 19294 22146 19346 22158
rect 15474 22094 15486 22146
rect 15538 22094 15550 22146
rect 15810 22094 15822 22146
rect 15874 22094 15886 22146
rect 13918 22082 13970 22094
rect 19294 22082 19346 22094
rect 23774 22146 23826 22158
rect 23774 22082 23826 22094
rect 24558 22146 24610 22158
rect 24558 22082 24610 22094
rect 27806 22146 27858 22158
rect 27806 22082 27858 22094
rect 28030 22146 28082 22158
rect 28030 22082 28082 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 15710 21810 15762 21822
rect 15362 21758 15374 21810
rect 15426 21758 15438 21810
rect 15710 21746 15762 21758
rect 17614 21810 17666 21822
rect 17614 21746 17666 21758
rect 17502 21698 17554 21710
rect 12114 21646 12126 21698
rect 12178 21646 12190 21698
rect 27906 21646 27918 21698
rect 27970 21646 27982 21698
rect 17502 21634 17554 21646
rect 18734 21586 18786 21598
rect 11330 21534 11342 21586
rect 11394 21534 11406 21586
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 18274 21534 18286 21586
rect 18338 21534 18350 21586
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 27122 21534 27134 21586
rect 27186 21534 27198 21586
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 18734 21522 18786 21534
rect 14702 21474 14754 21486
rect 14242 21422 14254 21474
rect 14306 21422 14318 21474
rect 14702 21410 14754 21422
rect 16830 21474 16882 21486
rect 23314 21422 23326 21474
rect 23378 21422 23390 21474
rect 30034 21422 30046 21474
rect 30098 21422 30110 21474
rect 16830 21410 16882 21422
rect 40014 21362 40066 21374
rect 40014 21298 40066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 22654 21026 22706 21038
rect 21970 20974 21982 21026
rect 22034 20974 22046 21026
rect 22654 20962 22706 20974
rect 15150 20914 15202 20926
rect 25330 20862 25342 20914
rect 25394 20862 25406 20914
rect 15150 20850 15202 20862
rect 21422 20802 21474 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 21422 20738 21474 20750
rect 21646 20802 21698 20814
rect 22642 20750 22654 20802
rect 22706 20750 22718 20802
rect 23314 20750 23326 20802
rect 23378 20750 23390 20802
rect 21646 20738 21698 20750
rect 22318 20690 22370 20702
rect 17490 20638 17502 20690
rect 17554 20638 17566 20690
rect 22318 20626 22370 20638
rect 14590 20578 14642 20590
rect 14590 20514 14642 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 17950 20242 18002 20254
rect 17950 20178 18002 20190
rect 22542 20242 22594 20254
rect 22542 20178 22594 20190
rect 14590 20130 14642 20142
rect 19854 20130 19906 20142
rect 15586 20078 15598 20130
rect 15650 20078 15662 20130
rect 14590 20066 14642 20078
rect 19854 20066 19906 20078
rect 21870 20130 21922 20142
rect 25230 20130 25282 20142
rect 23762 20078 23774 20130
rect 23826 20078 23838 20130
rect 21870 20066 21922 20078
rect 25230 20066 25282 20078
rect 15262 20018 15314 20030
rect 11330 19966 11342 20018
rect 11394 19966 11406 20018
rect 15262 19954 15314 19966
rect 16270 20018 16322 20030
rect 16270 19954 16322 19966
rect 18622 20018 18674 20030
rect 19282 19966 19294 20018
rect 19346 19966 19358 20018
rect 21298 19966 21310 20018
rect 21362 19966 21374 20018
rect 23538 19966 23550 20018
rect 23602 19966 23614 20018
rect 27458 19966 27470 20018
rect 27522 19966 27534 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 18622 19954 18674 19966
rect 16494 19906 16546 19918
rect 12002 19854 12014 19906
rect 12066 19854 12078 19906
rect 14130 19854 14142 19906
rect 14194 19854 14206 19906
rect 14466 19854 14478 19906
rect 14530 19854 14542 19906
rect 16494 19842 16546 19854
rect 17390 19906 17442 19918
rect 17390 19842 17442 19854
rect 25342 19906 25394 19918
rect 28242 19854 28254 19906
rect 28306 19854 28318 19906
rect 30370 19854 30382 19906
rect 30434 19854 30446 19906
rect 25342 19842 25394 19854
rect 14814 19794 14866 19806
rect 18734 19794 18786 19806
rect 15922 19742 15934 19794
rect 15986 19742 15998 19794
rect 14814 19730 14866 19742
rect 18734 19730 18786 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 21534 19458 21586 19470
rect 17938 19406 17950 19458
rect 18002 19406 18014 19458
rect 21534 19394 21586 19406
rect 21758 19458 21810 19470
rect 21758 19394 21810 19406
rect 14814 19346 14866 19358
rect 27470 19346 27522 19358
rect 22082 19294 22094 19346
rect 22146 19294 22158 19346
rect 23650 19294 23662 19346
rect 23714 19294 23726 19346
rect 25778 19294 25790 19346
rect 25842 19294 25854 19346
rect 14814 19282 14866 19294
rect 27470 19282 27522 19294
rect 40014 19346 40066 19358
rect 40014 19282 40066 19294
rect 14478 19234 14530 19246
rect 14478 19170 14530 19182
rect 16046 19234 16098 19246
rect 19070 19234 19122 19246
rect 22206 19234 22258 19246
rect 26686 19234 26738 19246
rect 17602 19182 17614 19234
rect 17666 19182 17678 19234
rect 19506 19182 19518 19234
rect 19570 19182 19582 19234
rect 22866 19182 22878 19234
rect 22930 19182 22942 19234
rect 16046 19170 16098 19182
rect 19070 19170 19122 19182
rect 22206 19170 22258 19182
rect 26686 19170 26738 19182
rect 27358 19234 27410 19246
rect 27358 19170 27410 19182
rect 27918 19234 27970 19246
rect 27918 19170 27970 19182
rect 28590 19234 28642 19246
rect 28590 19170 28642 19182
rect 29262 19234 29314 19246
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 29262 19170 29314 19182
rect 14590 19122 14642 19134
rect 14590 19058 14642 19070
rect 14926 19122 14978 19134
rect 14926 19058 14978 19070
rect 17054 19122 17106 19134
rect 22318 19122 22370 19134
rect 18162 19070 18174 19122
rect 18226 19070 18238 19122
rect 17054 19058 17106 19070
rect 22318 19058 22370 19070
rect 28366 19122 28418 19134
rect 28366 19058 28418 19070
rect 29374 19122 29426 19134
rect 29374 19058 29426 19070
rect 29710 19122 29762 19134
rect 29710 19058 29762 19070
rect 29934 19122 29986 19134
rect 29934 19058 29986 19070
rect 30158 19122 30210 19134
rect 30158 19058 30210 19070
rect 30270 19122 30322 19134
rect 30270 19058 30322 19070
rect 30606 19122 30658 19134
rect 30606 19058 30658 19070
rect 30718 19122 30770 19134
rect 30718 19058 30770 19070
rect 13806 19010 13858 19022
rect 13806 18946 13858 18958
rect 15374 19010 15426 19022
rect 16718 19010 16770 19022
rect 15698 18958 15710 19010
rect 15762 18958 15774 19010
rect 15374 18946 15426 18958
rect 16718 18946 16770 18958
rect 16942 19010 16994 19022
rect 16942 18946 16994 18958
rect 26910 19010 26962 19022
rect 26910 18946 26962 18958
rect 27134 19010 27186 19022
rect 27134 18946 27186 18958
rect 28254 19010 28306 19022
rect 28254 18946 28306 18958
rect 29486 19010 29538 19022
rect 29486 18946 29538 18958
rect 30942 19010 30994 19022
rect 30942 18946 30994 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 14030 18674 14082 18686
rect 26126 18674 26178 18686
rect 17826 18622 17838 18674
rect 17890 18622 17902 18674
rect 23650 18622 23662 18674
rect 23714 18622 23726 18674
rect 14030 18610 14082 18622
rect 26126 18610 26178 18622
rect 27358 18674 27410 18686
rect 27358 18610 27410 18622
rect 14254 18562 14306 18574
rect 25902 18562 25954 18574
rect 14578 18510 14590 18562
rect 14642 18510 14654 18562
rect 14254 18498 14306 18510
rect 25902 18498 25954 18510
rect 26350 18562 26402 18574
rect 26350 18498 26402 18510
rect 27022 18562 27074 18574
rect 27022 18498 27074 18510
rect 27134 18562 27186 18574
rect 28466 18510 28478 18562
rect 28530 18510 28542 18562
rect 27134 18498 27186 18510
rect 18174 18450 18226 18462
rect 22318 18450 22370 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 13570 18398 13582 18450
rect 13634 18398 13646 18450
rect 14466 18398 14478 18450
rect 14530 18398 14542 18450
rect 18610 18398 18622 18450
rect 18674 18398 18686 18450
rect 19394 18398 19406 18450
rect 19458 18398 19470 18450
rect 20402 18398 20414 18450
rect 20466 18398 20478 18450
rect 18174 18386 18226 18398
rect 22318 18386 22370 18398
rect 22654 18450 22706 18462
rect 22654 18386 22706 18398
rect 22990 18450 23042 18462
rect 22990 18386 23042 18398
rect 23326 18450 23378 18462
rect 23326 18386 23378 18398
rect 26462 18450 26514 18462
rect 27794 18398 27806 18450
rect 27858 18398 27870 18450
rect 26462 18386 26514 18398
rect 14142 18338 14194 18350
rect 10658 18286 10670 18338
rect 10722 18286 10734 18338
rect 12786 18286 12798 18338
rect 12850 18286 12862 18338
rect 14142 18274 14194 18286
rect 16494 18338 16546 18350
rect 17502 18338 17554 18350
rect 22542 18338 22594 18350
rect 16818 18286 16830 18338
rect 16882 18286 16894 18338
rect 18946 18286 18958 18338
rect 19010 18286 19022 18338
rect 20290 18286 20302 18338
rect 20354 18286 20366 18338
rect 30594 18286 30606 18338
rect 30658 18286 30670 18338
rect 16494 18274 16546 18286
rect 17502 18274 17554 18286
rect 22542 18274 22594 18286
rect 1934 18226 1986 18238
rect 20402 18174 20414 18226
rect 20466 18174 20478 18226
rect 1934 18162 1986 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 12462 17890 12514 17902
rect 12462 17826 12514 17838
rect 17054 17890 17106 17902
rect 17054 17826 17106 17838
rect 19294 17890 19346 17902
rect 19294 17826 19346 17838
rect 19518 17890 19570 17902
rect 19518 17826 19570 17838
rect 12350 17778 12402 17790
rect 16370 17726 16382 17778
rect 16434 17726 16446 17778
rect 22418 17726 22430 17778
rect 22482 17726 22494 17778
rect 24546 17726 24558 17778
rect 24610 17726 24622 17778
rect 12350 17714 12402 17726
rect 17726 17666 17778 17678
rect 13570 17614 13582 17666
rect 13634 17614 13646 17666
rect 17378 17614 17390 17666
rect 17442 17614 17454 17666
rect 19058 17614 19070 17666
rect 19122 17614 19134 17666
rect 21746 17614 21758 17666
rect 21810 17614 21822 17666
rect 17726 17602 17778 17614
rect 19630 17554 19682 17566
rect 14242 17502 14254 17554
rect 14306 17502 14318 17554
rect 18050 17502 18062 17554
rect 18114 17502 18126 17554
rect 19630 17490 19682 17502
rect 17166 17442 17218 17454
rect 17166 17378 17218 17390
rect 18398 17442 18450 17454
rect 18722 17390 18734 17442
rect 18786 17390 18798 17442
rect 18398 17378 18450 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 17838 17106 17890 17118
rect 17838 17042 17890 17054
rect 19854 17106 19906 17118
rect 22542 17106 22594 17118
rect 21410 17054 21422 17106
rect 21474 17054 21486 17106
rect 19854 17042 19906 17054
rect 22542 17042 22594 17054
rect 22654 17106 22706 17118
rect 22654 17042 22706 17054
rect 23438 17106 23490 17118
rect 23438 17042 23490 17054
rect 23662 17106 23714 17118
rect 23662 17042 23714 17054
rect 24222 17106 24274 17118
rect 24222 17042 24274 17054
rect 28366 17106 28418 17118
rect 28366 17042 28418 17054
rect 15038 16994 15090 17006
rect 15038 16930 15090 16942
rect 15262 16994 15314 17006
rect 20862 16994 20914 17006
rect 18274 16942 18286 16994
rect 18338 16942 18350 16994
rect 15262 16930 15314 16942
rect 20862 16930 20914 16942
rect 22206 16994 22258 17006
rect 22206 16930 22258 16942
rect 22766 16994 22818 17006
rect 26462 16994 26514 17006
rect 24546 16942 24558 16994
rect 24610 16942 24622 16994
rect 22766 16930 22818 16942
rect 26462 16930 26514 16942
rect 27358 16994 27410 17006
rect 27358 16930 27410 16942
rect 14926 16882 14978 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 14926 16818 14978 16830
rect 15486 16882 15538 16894
rect 17390 16882 17442 16894
rect 16818 16830 16830 16882
rect 16882 16830 16894 16882
rect 15486 16818 15538 16830
rect 17390 16818 17442 16830
rect 17614 16882 17666 16894
rect 22430 16882 22482 16894
rect 26686 16882 26738 16894
rect 28478 16882 28530 16894
rect 18498 16830 18510 16882
rect 18562 16830 18574 16882
rect 23202 16830 23214 16882
rect 23266 16830 23278 16882
rect 23874 16830 23886 16882
rect 23938 16830 23950 16882
rect 25778 16830 25790 16882
rect 25842 16830 25854 16882
rect 27122 16830 27134 16882
rect 27186 16830 27198 16882
rect 28018 16830 28030 16882
rect 28082 16830 28094 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 17614 16818 17666 16830
rect 22430 16818 22482 16830
rect 26686 16818 26738 16830
rect 28478 16818 28530 16830
rect 16606 16770 16658 16782
rect 16606 16706 16658 16718
rect 17502 16770 17554 16782
rect 17502 16706 17554 16718
rect 19630 16770 19682 16782
rect 19630 16706 19682 16718
rect 23550 16770 23602 16782
rect 23550 16706 23602 16718
rect 26014 16770 26066 16782
rect 26014 16706 26066 16718
rect 26574 16770 26626 16782
rect 26574 16706 26626 16718
rect 27694 16770 27746 16782
rect 27694 16706 27746 16718
rect 27806 16770 27858 16782
rect 39890 16718 39902 16770
rect 39954 16718 39966 16770
rect 27806 16706 27858 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 16494 16658 16546 16670
rect 16494 16594 16546 16606
rect 19966 16658 20018 16670
rect 19966 16594 20018 16606
rect 21086 16658 21138 16670
rect 21086 16594 21138 16606
rect 26126 16658 26178 16670
rect 26126 16594 26178 16606
rect 26910 16658 26962 16670
rect 26910 16594 26962 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 17838 16322 17890 16334
rect 17838 16258 17890 16270
rect 23438 16322 23490 16334
rect 23438 16258 23490 16270
rect 23774 16322 23826 16334
rect 23774 16258 23826 16270
rect 18062 16210 18114 16222
rect 23886 16210 23938 16222
rect 40014 16210 40066 16222
rect 23090 16158 23102 16210
rect 23154 16158 23166 16210
rect 26450 16158 26462 16210
rect 26514 16158 26526 16210
rect 28578 16158 28590 16210
rect 28642 16158 28654 16210
rect 18062 16146 18114 16158
rect 23886 16146 23938 16158
rect 40014 16146 40066 16158
rect 15822 16098 15874 16110
rect 15822 16034 15874 16046
rect 17278 16098 17330 16110
rect 25666 16046 25678 16098
rect 25730 16046 25742 16098
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 17278 16034 17330 16046
rect 15374 15986 15426 15998
rect 15374 15922 15426 15934
rect 15598 15986 15650 15998
rect 18286 15986 18338 15998
rect 17602 15934 17614 15986
rect 17666 15934 17678 15986
rect 15598 15922 15650 15934
rect 18286 15922 18338 15934
rect 23214 15986 23266 15998
rect 23214 15922 23266 15934
rect 15710 15874 15762 15886
rect 15710 15810 15762 15822
rect 18174 15874 18226 15886
rect 18174 15810 18226 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 18510 15538 18562 15550
rect 18510 15474 18562 15486
rect 16270 15426 16322 15438
rect 20638 15426 20690 15438
rect 19282 15374 19294 15426
rect 19346 15374 19358 15426
rect 16270 15362 16322 15374
rect 20638 15362 20690 15374
rect 20750 15426 20802 15438
rect 22530 15374 22542 15426
rect 22594 15374 22606 15426
rect 26002 15374 26014 15426
rect 26066 15374 26078 15426
rect 20750 15362 20802 15374
rect 16046 15314 16098 15326
rect 15362 15262 15374 15314
rect 15426 15262 15438 15314
rect 16046 15250 16098 15262
rect 18622 15314 18674 15326
rect 18622 15250 18674 15262
rect 18958 15314 19010 15326
rect 18958 15250 19010 15262
rect 19742 15314 19794 15326
rect 19742 15250 19794 15262
rect 19966 15314 20018 15326
rect 20178 15262 20190 15314
rect 20242 15262 20254 15314
rect 21858 15262 21870 15314
rect 21922 15262 21934 15314
rect 25330 15262 25342 15314
rect 25394 15262 25406 15314
rect 19966 15250 20018 15262
rect 15710 15202 15762 15214
rect 12450 15150 12462 15202
rect 12514 15150 12526 15202
rect 14578 15150 14590 15202
rect 14642 15150 14654 15202
rect 15710 15138 15762 15150
rect 20526 15202 20578 15214
rect 24658 15150 24670 15202
rect 24722 15150 24734 15202
rect 28130 15150 28142 15202
rect 28194 15150 28206 15202
rect 20526 15138 20578 15150
rect 19630 15090 19682 15102
rect 19630 15026 19682 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 14142 14754 14194 14766
rect 14142 14690 14194 14702
rect 14030 14642 14082 14654
rect 20738 14590 20750 14642
rect 20802 14590 20814 14642
rect 14030 14578 14082 14590
rect 17826 14478 17838 14530
rect 17890 14478 17902 14530
rect 18610 14478 18622 14530
rect 18674 14478 18686 14530
rect 15598 14306 15650 14318
rect 15598 14242 15650 14254
rect 17502 14306 17554 14318
rect 17502 14242 17554 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 18162 13806 18174 13858
rect 18226 13806 18238 13858
rect 20750 13746 20802 13758
rect 17490 13694 17502 13746
rect 17554 13694 17566 13746
rect 20750 13682 20802 13694
rect 20290 13582 20302 13634
rect 20354 13582 20366 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 24782 5234 24834 5246
rect 24782 5170 24834 5182
rect 23762 5070 23774 5122
rect 23826 5070 23838 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 19730 4286 19742 4338
rect 19794 4286 19806 4338
rect 20750 4114 20802 4126
rect 20750 4050 20802 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 18834 3614 18846 3666
rect 18898 3614 18910 3666
rect 25566 3602 25618 3614
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 35982 3330 36034 3342
rect 35982 3266 36034 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 26126 38222 26178 38274
rect 18846 38110 18898 38162
rect 22206 38110 22258 38162
rect 17614 37998 17666 38050
rect 23550 37998 23602 38050
rect 25566 37998 25618 38050
rect 30494 37886 30546 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 22766 37438 22818 37490
rect 26798 37438 26850 37490
rect 20974 37214 21026 37266
rect 22206 37214 22258 37266
rect 25902 37214 25954 37266
rect 19518 37102 19570 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 16718 36654 16770 36706
rect 15710 36430 15762 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 22542 28030 22594 28082
rect 22878 28030 22930 28082
rect 23774 27918 23826 27970
rect 19294 27806 19346 27858
rect 23662 27806 23714 27858
rect 17838 27694 17890 27746
rect 19070 27694 19122 27746
rect 20078 27694 20130 27746
rect 22206 27694 22258 27746
rect 17726 27582 17778 27634
rect 23774 27582 23826 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1934 27134 1986 27186
rect 16942 27134 16994 27186
rect 19070 27134 19122 27186
rect 23774 27134 23826 27186
rect 25902 27134 25954 27186
rect 4286 27022 4338 27074
rect 16158 27022 16210 27074
rect 22990 27022 23042 27074
rect 14254 26910 14306 26962
rect 14366 26910 14418 26962
rect 19518 26910 19570 26962
rect 19630 26910 19682 26962
rect 19294 26798 19346 26850
rect 20078 26798 20130 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 20862 26462 20914 26514
rect 21422 26462 21474 26514
rect 23886 26462 23938 26514
rect 24558 26462 24610 26514
rect 13358 26350 13410 26402
rect 20750 26350 20802 26402
rect 12686 26238 12738 26290
rect 15934 26238 15986 26290
rect 16046 26238 16098 26290
rect 16158 26238 16210 26290
rect 16270 26238 16322 26290
rect 16382 26238 16434 26290
rect 17390 26238 17442 26290
rect 23438 26238 23490 26290
rect 23662 26238 23714 26290
rect 23998 26238 24050 26290
rect 24446 26238 24498 26290
rect 15486 26126 15538 26178
rect 18174 26126 18226 26178
rect 20302 26126 20354 26178
rect 22990 26126 23042 26178
rect 23774 26126 23826 26178
rect 20862 26014 20914 26066
rect 23102 26014 23154 26066
rect 24558 26014 24610 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 15486 25678 15538 25730
rect 15934 25678 15986 25730
rect 19406 25678 19458 25730
rect 22430 25678 22482 25730
rect 13470 25566 13522 25618
rect 14590 25566 14642 25618
rect 16270 25566 16322 25618
rect 20190 25566 20242 25618
rect 23662 25566 23714 25618
rect 25790 25566 25842 25618
rect 14702 25454 14754 25506
rect 17502 25454 17554 25506
rect 17726 25454 17778 25506
rect 17950 25454 18002 25506
rect 18174 25454 18226 25506
rect 18622 25454 18674 25506
rect 18846 25454 18898 25506
rect 19854 25454 19906 25506
rect 20638 25454 20690 25506
rect 22878 25454 22930 25506
rect 15150 25342 15202 25394
rect 16270 25342 16322 25394
rect 16494 25342 16546 25394
rect 17278 25342 17330 25394
rect 19182 25342 19234 25394
rect 20078 25342 20130 25394
rect 20190 25342 20242 25394
rect 22430 25342 22482 25394
rect 22542 25342 22594 25394
rect 13582 25230 13634 25282
rect 14590 25230 14642 25282
rect 14926 25230 14978 25282
rect 15710 25230 15762 25282
rect 17726 25230 17778 25282
rect 18510 25230 18562 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 20414 24894 20466 24946
rect 22654 24894 22706 24946
rect 13918 24782 13970 24834
rect 18398 24782 18450 24834
rect 14590 24670 14642 24722
rect 15150 24670 15202 24722
rect 18734 24670 18786 24722
rect 18958 24670 19010 24722
rect 20750 24670 20802 24722
rect 22318 24670 22370 24722
rect 26574 24670 26626 24722
rect 37662 24670 37714 24722
rect 11790 24558 11842 24610
rect 27358 24558 27410 24610
rect 29486 24558 29538 24610
rect 18510 24446 18562 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 27470 24110 27522 24162
rect 40014 23998 40066 24050
rect 37662 23886 37714 23938
rect 18510 23774 18562 23826
rect 19294 23774 19346 23826
rect 22654 23774 22706 23826
rect 27582 23774 27634 23826
rect 28030 23774 28082 23826
rect 28254 23774 28306 23826
rect 28366 23774 28418 23826
rect 14366 23662 14418 23714
rect 18622 23662 18674 23714
rect 18958 23662 19010 23714
rect 22542 23662 22594 23714
rect 27470 23662 27522 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 19630 23326 19682 23378
rect 20862 23326 20914 23378
rect 12014 23214 12066 23266
rect 17390 23214 17442 23266
rect 19182 23214 19234 23266
rect 19966 23214 20018 23266
rect 11342 23102 11394 23154
rect 14926 23102 14978 23154
rect 17726 23102 17778 23154
rect 18174 23102 18226 23154
rect 19070 23102 19122 23154
rect 20638 23102 20690 23154
rect 21870 23102 21922 23154
rect 27134 23102 27186 23154
rect 37662 23102 37714 23154
rect 14142 22990 14194 23042
rect 14478 22990 14530 23042
rect 15374 22990 15426 23042
rect 18622 22990 18674 23042
rect 22542 22990 22594 23042
rect 24670 22990 24722 23042
rect 27918 22990 27970 23042
rect 30046 22990 30098 23042
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 15150 22542 15202 22594
rect 28478 22542 28530 22594
rect 16382 22430 16434 22482
rect 18958 22430 19010 22482
rect 21310 22430 21362 22482
rect 28590 22430 28642 22482
rect 29262 22430 29314 22482
rect 40014 22430 40066 22482
rect 14254 22318 14306 22370
rect 14926 22318 14978 22370
rect 16158 22318 16210 22370
rect 17390 22318 17442 22370
rect 19182 22318 19234 22370
rect 22318 22318 22370 22370
rect 23438 22318 23490 22370
rect 23662 22318 23714 22370
rect 24446 22318 24498 22370
rect 27694 22318 27746 22370
rect 28142 22318 28194 22370
rect 29038 22318 29090 22370
rect 29486 22318 29538 22370
rect 29598 22318 29650 22370
rect 37662 22318 37714 22370
rect 17838 22206 17890 22258
rect 20190 22206 20242 22258
rect 21646 22206 21698 22258
rect 22654 22206 22706 22258
rect 22990 22206 23042 22258
rect 23214 22206 23266 22258
rect 23886 22206 23938 22258
rect 24222 22206 24274 22258
rect 24782 22206 24834 22258
rect 27358 22206 27410 22258
rect 27470 22206 27522 22258
rect 13918 22094 13970 22146
rect 15486 22094 15538 22146
rect 15822 22094 15874 22146
rect 19294 22094 19346 22146
rect 23774 22094 23826 22146
rect 24558 22094 24610 22146
rect 27806 22094 27858 22146
rect 28030 22094 28082 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 15374 21758 15426 21810
rect 15710 21758 15762 21810
rect 17614 21758 17666 21810
rect 12126 21646 12178 21698
rect 17502 21646 17554 21698
rect 27918 21646 27970 21698
rect 11342 21534 11394 21586
rect 17838 21534 17890 21586
rect 18286 21534 18338 21586
rect 18734 21534 18786 21586
rect 19406 21534 19458 21586
rect 27134 21534 27186 21586
rect 37886 21534 37938 21586
rect 14254 21422 14306 21474
rect 14702 21422 14754 21474
rect 16830 21422 16882 21474
rect 23326 21422 23378 21474
rect 30046 21422 30098 21474
rect 40014 21310 40066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 21982 20974 22034 21026
rect 22654 20974 22706 21026
rect 15150 20862 15202 20914
rect 25342 20862 25394 20914
rect 20078 20750 20130 20802
rect 21422 20750 21474 20802
rect 21646 20750 21698 20802
rect 22654 20750 22706 20802
rect 23326 20750 23378 20802
rect 17502 20638 17554 20690
rect 22318 20638 22370 20690
rect 14590 20526 14642 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 17950 20190 18002 20242
rect 22542 20190 22594 20242
rect 14590 20078 14642 20130
rect 15598 20078 15650 20130
rect 19854 20078 19906 20130
rect 21870 20078 21922 20130
rect 23774 20078 23826 20130
rect 25230 20078 25282 20130
rect 11342 19966 11394 20018
rect 15262 19966 15314 20018
rect 16270 19966 16322 20018
rect 18622 19966 18674 20018
rect 19294 19966 19346 20018
rect 21310 19966 21362 20018
rect 23550 19966 23602 20018
rect 27470 19966 27522 20018
rect 37662 19966 37714 20018
rect 12014 19854 12066 19906
rect 14142 19854 14194 19906
rect 14478 19854 14530 19906
rect 16494 19854 16546 19906
rect 17390 19854 17442 19906
rect 25342 19854 25394 19906
rect 28254 19854 28306 19906
rect 30382 19854 30434 19906
rect 14814 19742 14866 19794
rect 15934 19742 15986 19794
rect 18734 19742 18786 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 17950 19406 18002 19458
rect 21534 19406 21586 19458
rect 21758 19406 21810 19458
rect 14814 19294 14866 19346
rect 22094 19294 22146 19346
rect 23662 19294 23714 19346
rect 25790 19294 25842 19346
rect 27470 19294 27522 19346
rect 40014 19294 40066 19346
rect 14478 19182 14530 19234
rect 16046 19182 16098 19234
rect 17614 19182 17666 19234
rect 19070 19182 19122 19234
rect 19518 19182 19570 19234
rect 22206 19182 22258 19234
rect 22878 19182 22930 19234
rect 26686 19182 26738 19234
rect 27358 19182 27410 19234
rect 27918 19182 27970 19234
rect 28590 19182 28642 19234
rect 29262 19182 29314 19234
rect 37662 19182 37714 19234
rect 14590 19070 14642 19122
rect 14926 19070 14978 19122
rect 17054 19070 17106 19122
rect 18174 19070 18226 19122
rect 22318 19070 22370 19122
rect 28366 19070 28418 19122
rect 29374 19070 29426 19122
rect 29710 19070 29762 19122
rect 29934 19070 29986 19122
rect 30158 19070 30210 19122
rect 30270 19070 30322 19122
rect 30606 19070 30658 19122
rect 30718 19070 30770 19122
rect 13806 18958 13858 19010
rect 15374 18958 15426 19010
rect 15710 18958 15762 19010
rect 16718 18958 16770 19010
rect 16942 18958 16994 19010
rect 26910 18958 26962 19010
rect 27134 18958 27186 19010
rect 28254 18958 28306 19010
rect 29486 18958 29538 19010
rect 30942 18958 30994 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 14030 18622 14082 18674
rect 17838 18622 17890 18674
rect 23662 18622 23714 18674
rect 26126 18622 26178 18674
rect 27358 18622 27410 18674
rect 14254 18510 14306 18562
rect 14590 18510 14642 18562
rect 25902 18510 25954 18562
rect 26350 18510 26402 18562
rect 27022 18510 27074 18562
rect 27134 18510 27186 18562
rect 28478 18510 28530 18562
rect 4286 18398 4338 18450
rect 13582 18398 13634 18450
rect 14478 18398 14530 18450
rect 18174 18398 18226 18450
rect 18622 18398 18674 18450
rect 19406 18398 19458 18450
rect 20414 18398 20466 18450
rect 22318 18398 22370 18450
rect 22654 18398 22706 18450
rect 22990 18398 23042 18450
rect 23326 18398 23378 18450
rect 26462 18398 26514 18450
rect 27806 18398 27858 18450
rect 10670 18286 10722 18338
rect 12798 18286 12850 18338
rect 14142 18286 14194 18338
rect 16494 18286 16546 18338
rect 16830 18286 16882 18338
rect 17502 18286 17554 18338
rect 18958 18286 19010 18338
rect 20302 18286 20354 18338
rect 22542 18286 22594 18338
rect 30606 18286 30658 18338
rect 1934 18174 1986 18226
rect 20414 18174 20466 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 12462 17838 12514 17890
rect 17054 17838 17106 17890
rect 19294 17838 19346 17890
rect 19518 17838 19570 17890
rect 12350 17726 12402 17778
rect 16382 17726 16434 17778
rect 22430 17726 22482 17778
rect 24558 17726 24610 17778
rect 13582 17614 13634 17666
rect 17390 17614 17442 17666
rect 17726 17614 17778 17666
rect 19070 17614 19122 17666
rect 21758 17614 21810 17666
rect 14254 17502 14306 17554
rect 18062 17502 18114 17554
rect 19630 17502 19682 17554
rect 17166 17390 17218 17442
rect 18398 17390 18450 17442
rect 18734 17390 18786 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17838 17054 17890 17106
rect 19854 17054 19906 17106
rect 21422 17054 21474 17106
rect 22542 17054 22594 17106
rect 22654 17054 22706 17106
rect 23438 17054 23490 17106
rect 23662 17054 23714 17106
rect 24222 17054 24274 17106
rect 28366 17054 28418 17106
rect 15038 16942 15090 16994
rect 15262 16942 15314 16994
rect 18286 16942 18338 16994
rect 20862 16942 20914 16994
rect 22206 16942 22258 16994
rect 22766 16942 22818 16994
rect 24558 16942 24610 16994
rect 26462 16942 26514 16994
rect 27358 16942 27410 16994
rect 4286 16830 4338 16882
rect 14926 16830 14978 16882
rect 15486 16830 15538 16882
rect 16830 16830 16882 16882
rect 17390 16830 17442 16882
rect 17614 16830 17666 16882
rect 18510 16830 18562 16882
rect 22430 16830 22482 16882
rect 23214 16830 23266 16882
rect 23886 16830 23938 16882
rect 25790 16830 25842 16882
rect 26686 16830 26738 16882
rect 27134 16830 27186 16882
rect 28030 16830 28082 16882
rect 28478 16830 28530 16882
rect 37662 16830 37714 16882
rect 16606 16718 16658 16770
rect 17502 16718 17554 16770
rect 19630 16718 19682 16770
rect 23550 16718 23602 16770
rect 26014 16718 26066 16770
rect 26574 16718 26626 16770
rect 27694 16718 27746 16770
rect 27806 16718 27858 16770
rect 39902 16718 39954 16770
rect 1934 16606 1986 16658
rect 16494 16606 16546 16658
rect 19966 16606 20018 16658
rect 21086 16606 21138 16658
rect 26126 16606 26178 16658
rect 26910 16606 26962 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 17838 16270 17890 16322
rect 23438 16270 23490 16322
rect 23774 16270 23826 16322
rect 18062 16158 18114 16210
rect 23102 16158 23154 16210
rect 23886 16158 23938 16210
rect 26462 16158 26514 16210
rect 28590 16158 28642 16210
rect 40014 16158 40066 16210
rect 15822 16046 15874 16098
rect 17278 16046 17330 16098
rect 25678 16046 25730 16098
rect 37662 16046 37714 16098
rect 15374 15934 15426 15986
rect 15598 15934 15650 15986
rect 17614 15934 17666 15986
rect 18286 15934 18338 15986
rect 23214 15934 23266 15986
rect 15710 15822 15762 15874
rect 18174 15822 18226 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 18510 15486 18562 15538
rect 16270 15374 16322 15426
rect 19294 15374 19346 15426
rect 20638 15374 20690 15426
rect 20750 15374 20802 15426
rect 22542 15374 22594 15426
rect 26014 15374 26066 15426
rect 15374 15262 15426 15314
rect 16046 15262 16098 15314
rect 18622 15262 18674 15314
rect 18958 15262 19010 15314
rect 19742 15262 19794 15314
rect 19966 15262 20018 15314
rect 20190 15262 20242 15314
rect 21870 15262 21922 15314
rect 25342 15262 25394 15314
rect 12462 15150 12514 15202
rect 14590 15150 14642 15202
rect 15710 15150 15762 15202
rect 20526 15150 20578 15202
rect 24670 15150 24722 15202
rect 28142 15150 28194 15202
rect 19630 15038 19682 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 14142 14702 14194 14754
rect 14030 14590 14082 14642
rect 20750 14590 20802 14642
rect 17838 14478 17890 14530
rect 18622 14478 18674 14530
rect 15598 14254 15650 14306
rect 17502 14254 17554 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 18174 13806 18226 13858
rect 17502 13694 17554 13746
rect 20750 13694 20802 13746
rect 20302 13582 20354 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 24782 5182 24834 5234
rect 23774 5070 23826 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19742 4286 19794 4338
rect 20750 4062 20802 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18846 3614 18898 3666
rect 25566 3614 25618 3666
rect 19742 3502 19794 3554
rect 20750 3502 20802 3554
rect 24558 3502 24610 3554
rect 21758 3278 21810 3330
rect 35982 3278 36034 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 15456 41200 15568 42000
rect 18816 41200 18928 42000
rect 19488 41200 19600 42000
rect 21504 41200 21616 42000
rect 22176 41200 22288 42000
rect 24864 41200 24976 42000
rect 25536 41200 25648 42000
rect 30240 41200 30352 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 15484 36708 15540 41200
rect 18844 38162 18900 41200
rect 18844 38110 18846 38162
rect 18898 38110 18900 38162
rect 18844 38098 18900 38110
rect 17612 38050 17668 38062
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 15484 36642 15540 36652
rect 16716 36708 16772 36718
rect 16716 36614 16772 36652
rect 15708 36482 15764 36494
rect 15708 36430 15710 36482
rect 15762 36430 15764 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 15708 31948 15764 36430
rect 15484 31892 15764 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4172 27636 4228 27646
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 1932 26226 1988 26236
rect 4172 21476 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 11788 27076 11844 27086
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 11788 25508 11844 27020
rect 13356 26964 13412 26974
rect 13356 26402 13412 26908
rect 14252 26964 14308 26974
rect 14252 26870 14308 26908
rect 14364 26962 14420 26974
rect 14364 26910 14366 26962
rect 14418 26910 14420 26962
rect 13356 26350 13358 26402
rect 13410 26350 13412 26402
rect 13356 26338 13412 26350
rect 11788 24610 11844 25452
rect 12684 26290 12740 26302
rect 12684 26238 12686 26290
rect 12738 26238 12740 26290
rect 12684 24724 12740 26238
rect 14364 26292 14420 26910
rect 14364 26226 14420 26236
rect 15484 26178 15540 31892
rect 17612 27860 17668 37998
rect 19516 37154 19572 41200
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 21532 37492 21588 41200
rect 22204 38162 22260 41200
rect 24892 38276 24948 41200
rect 25564 38612 25620 41200
rect 25564 38546 25620 38556
rect 26796 38612 26852 38622
rect 24892 38210 24948 38220
rect 26124 38276 26180 38286
rect 26124 38182 26180 38220
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 23548 38050 23604 38062
rect 23548 37998 23550 38050
rect 23602 37998 23604 38050
rect 21532 37426 21588 37436
rect 22764 37492 22820 37502
rect 22764 37398 22820 37436
rect 19516 37102 19518 37154
rect 19570 37102 19572 37154
rect 19516 37090 19572 37102
rect 20972 37266 21028 37278
rect 20972 37214 20974 37266
rect 21026 37214 21028 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 28532 19572 28542
rect 18172 27860 18228 27870
rect 17612 27794 17668 27804
rect 18060 27804 18172 27860
rect 17836 27746 17892 27758
rect 17836 27694 17838 27746
rect 17890 27694 17892 27746
rect 17724 27636 17780 27646
rect 16940 27634 17780 27636
rect 16940 27582 17726 27634
rect 17778 27582 17780 27634
rect 16940 27580 17780 27582
rect 16940 27186 16996 27580
rect 17724 27570 17780 27580
rect 16940 27134 16942 27186
rect 16994 27134 16996 27186
rect 16940 27122 16996 27134
rect 16156 27076 16212 27086
rect 15484 26126 15486 26178
rect 15538 26126 15540 26178
rect 14924 25956 14980 25966
rect 14812 25900 14924 25956
rect 13468 25620 13524 25630
rect 14588 25620 14644 25630
rect 13468 25618 14644 25620
rect 13468 25566 13470 25618
rect 13522 25566 14590 25618
rect 14642 25566 14644 25618
rect 13468 25564 14644 25566
rect 13468 25554 13524 25564
rect 14588 25554 14644 25564
rect 14700 25508 14756 25518
rect 14700 25414 14756 25452
rect 13580 25284 13636 25294
rect 14588 25284 14644 25294
rect 14812 25284 14868 25900
rect 14924 25890 14980 25900
rect 15484 25730 15540 26126
rect 15484 25678 15486 25730
rect 15538 25678 15540 25730
rect 15484 25666 15540 25678
rect 15820 27074 16212 27076
rect 15820 27022 16158 27074
rect 16210 27022 16212 27074
rect 15820 27020 16212 27022
rect 15820 26180 15876 27020
rect 16156 27010 16212 27020
rect 17388 26964 17444 26974
rect 15148 25394 15204 25406
rect 15148 25342 15150 25394
rect 15202 25342 15204 25394
rect 13580 25282 13972 25284
rect 13580 25230 13582 25282
rect 13634 25230 13972 25282
rect 13580 25228 13972 25230
rect 13580 25218 13636 25228
rect 13916 24834 13972 25228
rect 14588 25282 14868 25284
rect 14588 25230 14590 25282
rect 14642 25230 14868 25282
rect 14588 25228 14868 25230
rect 14924 25284 14980 25294
rect 15148 25284 15204 25342
rect 15372 25284 15428 25294
rect 14924 25282 15092 25284
rect 14924 25230 14926 25282
rect 14978 25230 15092 25282
rect 14924 25228 15092 25230
rect 15148 25228 15372 25284
rect 14588 25218 14644 25228
rect 14924 25218 14980 25228
rect 13916 24782 13918 24834
rect 13970 24782 13972 24834
rect 13916 24770 13972 24782
rect 12684 24658 12740 24668
rect 14588 24724 14644 24734
rect 11788 24558 11790 24610
rect 11842 24558 11844 24610
rect 11788 24546 11844 24558
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 14364 23714 14420 23726
rect 14364 23662 14366 23714
rect 14418 23662 14420 23714
rect 14364 23604 14420 23662
rect 14588 23604 14644 24668
rect 14364 23548 14644 23604
rect 12012 23380 12068 23390
rect 12012 23266 12068 23324
rect 12012 23214 12014 23266
rect 12066 23214 12068 23266
rect 12012 23202 12068 23214
rect 11340 23154 11396 23166
rect 11340 23102 11342 23154
rect 11394 23102 11396 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 21410 4228 21420
rect 11340 21586 11396 23102
rect 14140 23042 14196 23054
rect 14476 23044 14532 23054
rect 14140 22990 14142 23042
rect 14194 22990 14196 23042
rect 14140 22596 14196 22990
rect 14140 22530 14196 22540
rect 14252 23042 14532 23044
rect 14252 22990 14478 23042
rect 14530 22990 14532 23042
rect 14252 22988 14532 22990
rect 14140 22372 14196 22382
rect 12124 22148 12180 22158
rect 12124 21698 12180 22092
rect 13916 22148 13972 22158
rect 13916 22054 13972 22092
rect 12124 21646 12126 21698
rect 12178 21646 12180 21698
rect 12124 21634 12180 21646
rect 11340 21534 11342 21586
rect 11394 21534 11396 21586
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 11340 20018 11396 21534
rect 14140 21476 14196 22316
rect 14252 22370 14308 22988
rect 14476 22978 14532 22988
rect 14252 22318 14254 22370
rect 14306 22318 14308 22370
rect 14252 22306 14308 22318
rect 14252 21476 14308 21486
rect 14140 21474 14308 21476
rect 14140 21422 14254 21474
rect 14306 21422 14308 21474
rect 14140 21420 14308 21422
rect 14588 21476 14644 23548
rect 14924 23154 14980 23166
rect 14924 23102 14926 23154
rect 14978 23102 14980 23154
rect 14924 22596 14980 23102
rect 14924 22530 14980 22540
rect 14924 22370 14980 22382
rect 14924 22318 14926 22370
rect 14978 22318 14980 22370
rect 14924 22148 14980 22318
rect 14924 22082 14980 22092
rect 15036 21812 15092 25228
rect 15148 24724 15204 24762
rect 15148 24658 15204 24668
rect 15372 23492 15428 25228
rect 15708 25284 15764 25294
rect 15820 25284 15876 26124
rect 15932 26290 15988 26302
rect 15932 26238 15934 26290
rect 15986 26238 15988 26290
rect 15932 25956 15988 26238
rect 15932 25890 15988 25900
rect 16044 26290 16100 26302
rect 16044 26238 16046 26290
rect 16098 26238 16100 26290
rect 15932 25732 15988 25742
rect 16044 25732 16100 26238
rect 16156 26292 16212 26302
rect 16156 26198 16212 26236
rect 16268 26290 16324 26302
rect 16268 26238 16270 26290
rect 16322 26238 16324 26290
rect 15932 25730 16100 25732
rect 15932 25678 15934 25730
rect 15986 25678 16100 25730
rect 15932 25676 16100 25678
rect 15932 25666 15988 25676
rect 16268 25618 16324 26238
rect 16268 25566 16270 25618
rect 16322 25566 16324 25618
rect 16268 25554 16324 25566
rect 16380 26290 16436 26302
rect 16380 26238 16382 26290
rect 16434 26238 16436 26290
rect 16380 25508 16436 26238
rect 17388 26290 17444 26908
rect 17388 26238 17390 26290
rect 17442 26238 17444 26290
rect 17388 26180 17444 26238
rect 17388 26114 17444 26124
rect 16268 25396 16324 25406
rect 16268 25302 16324 25340
rect 15708 25282 15876 25284
rect 15708 25230 15710 25282
rect 15762 25230 15876 25282
rect 15708 25228 15876 25230
rect 16380 25284 16436 25452
rect 17500 25508 17556 25518
rect 17724 25508 17780 25518
rect 17500 25414 17556 25452
rect 17612 25506 17780 25508
rect 17612 25454 17726 25506
rect 17778 25454 17780 25506
rect 17612 25452 17780 25454
rect 15708 24724 15764 25228
rect 16380 25218 16436 25228
rect 16492 25394 16548 25406
rect 16492 25342 16494 25394
rect 16546 25342 16548 25394
rect 15708 24658 15764 24668
rect 16492 24724 16548 25342
rect 17276 25394 17332 25406
rect 17276 25342 17278 25394
rect 17330 25342 17332 25394
rect 17276 25284 17332 25342
rect 17276 25218 17332 25228
rect 17612 25060 17668 25452
rect 17724 25442 17780 25452
rect 17724 25284 17780 25294
rect 17836 25284 17892 27694
rect 17948 25508 18004 25518
rect 18060 25508 18116 27804
rect 18172 27794 18228 27804
rect 19292 27858 19348 27870
rect 19292 27806 19294 27858
rect 19346 27806 19348 27858
rect 19068 27748 19124 27758
rect 19292 27748 19348 27806
rect 18956 27746 19348 27748
rect 18956 27694 19070 27746
rect 19122 27694 19348 27746
rect 18956 27692 19348 27694
rect 18844 26964 18900 26974
rect 18956 26964 19012 27692
rect 19068 27682 19124 27692
rect 19068 27524 19124 27534
rect 19068 27186 19124 27468
rect 19068 27134 19070 27186
rect 19122 27134 19124 27186
rect 19068 27122 19124 27134
rect 18900 26908 19012 26964
rect 19516 27076 19572 28476
rect 20972 28532 21028 37214
rect 22204 37266 22260 37278
rect 22204 37214 22206 37266
rect 22258 37214 22260 37266
rect 22204 31948 22260 37214
rect 22204 31892 22932 31948
rect 20972 28466 21028 28476
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 22540 28084 22596 28094
rect 22876 28084 22932 31892
rect 22540 27990 22596 28028
rect 22652 28082 22932 28084
rect 22652 28030 22878 28082
rect 22930 28030 22932 28082
rect 22652 28028 22932 28030
rect 20076 27746 20132 27758
rect 20076 27694 20078 27746
rect 20130 27694 20132 27746
rect 20076 27076 20132 27694
rect 22204 27748 22260 27758
rect 22652 27748 22708 28028
rect 22876 28018 22932 28028
rect 23548 28084 23604 37998
rect 25564 38050 25620 38062
rect 25564 37998 25566 38050
rect 25618 37998 25620 38050
rect 25564 31948 25620 37998
rect 26796 37490 26852 38556
rect 30268 37940 30324 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 30492 37940 30548 37950
rect 30268 37938 30548 37940
rect 30268 37886 30494 37938
rect 30546 37886 30548 37938
rect 30268 37884 30548 37886
rect 30492 37874 30548 37884
rect 26796 37438 26798 37490
rect 26850 37438 26852 37490
rect 26796 37426 26852 37438
rect 25900 37266 25956 37278
rect 25900 37214 25902 37266
rect 25954 37214 25956 37266
rect 25564 31892 25844 31948
rect 23548 28018 23604 28028
rect 23772 27972 23828 27982
rect 23772 27970 24388 27972
rect 23772 27918 23774 27970
rect 23826 27918 24388 27970
rect 23772 27916 24388 27918
rect 23772 27906 23828 27916
rect 22204 27746 22708 27748
rect 22204 27694 22206 27746
rect 22258 27694 22708 27746
rect 22204 27692 22708 27694
rect 23660 27858 23716 27870
rect 23660 27806 23662 27858
rect 23714 27806 23716 27858
rect 20076 27020 20468 27076
rect 19516 26962 19572 27020
rect 19516 26910 19518 26962
rect 19570 26910 19572 26962
rect 18844 26898 18900 26908
rect 19516 26898 19572 26910
rect 19628 26962 19684 26974
rect 19628 26910 19630 26962
rect 19682 26910 19684 26962
rect 19292 26850 19348 26862
rect 19292 26798 19294 26850
rect 19346 26798 19348 26850
rect 18172 26180 18228 26190
rect 18172 26178 18340 26180
rect 18172 26126 18174 26178
rect 18226 26126 18340 26178
rect 18172 26124 18340 26126
rect 18172 26114 18228 26124
rect 18172 25508 18228 25518
rect 18060 25506 18228 25508
rect 18060 25454 18174 25506
rect 18226 25454 18228 25506
rect 18060 25452 18228 25454
rect 17948 25414 18004 25452
rect 18172 25442 18228 25452
rect 17724 25282 17892 25284
rect 17724 25230 17726 25282
rect 17778 25230 17892 25282
rect 17724 25228 17892 25230
rect 18284 25284 18340 26124
rect 19292 25732 19348 26798
rect 19628 26404 19684 26910
rect 19964 26964 20020 26974
rect 20020 26908 20132 26964
rect 19964 26898 20020 26908
rect 20076 26852 20132 26908
rect 20300 26852 20356 26862
rect 20076 26850 20244 26852
rect 20076 26798 20078 26850
rect 20130 26798 20244 26850
rect 20076 26796 20244 26798
rect 20076 26786 20132 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20188 26516 20244 26796
rect 20188 26450 20244 26460
rect 19628 26338 19684 26348
rect 20300 26178 20356 26796
rect 20300 26126 20302 26178
rect 20354 26126 20356 26178
rect 20300 26114 20356 26126
rect 19404 25732 19460 25742
rect 18620 25676 19236 25732
rect 19292 25730 19460 25732
rect 19292 25678 19406 25730
rect 19458 25678 19460 25730
rect 19292 25676 19460 25678
rect 18620 25506 18676 25676
rect 19180 25620 19236 25676
rect 19404 25666 19460 25676
rect 20188 25620 20244 25630
rect 20412 25620 20468 27020
rect 20860 26852 20916 26862
rect 20860 26514 20916 26796
rect 22204 26852 22260 27692
rect 22988 27076 23044 27086
rect 22876 27074 23044 27076
rect 22876 27022 22990 27074
rect 23042 27022 23044 27074
rect 22876 27020 23044 27022
rect 22204 26786 22260 26796
rect 22428 26964 22484 26974
rect 20860 26462 20862 26514
rect 20914 26462 20916 26514
rect 20860 26450 20916 26462
rect 21420 26516 21476 26526
rect 21420 26422 21476 26460
rect 19180 25564 19348 25620
rect 18620 25454 18622 25506
rect 18674 25454 18676 25506
rect 18508 25284 18564 25294
rect 18284 25282 18564 25284
rect 18284 25230 18510 25282
rect 18562 25230 18564 25282
rect 18284 25228 18564 25230
rect 17724 25218 17780 25228
rect 18508 25218 18564 25228
rect 17612 25004 18452 25060
rect 18396 24834 18452 25004
rect 18396 24782 18398 24834
rect 18450 24782 18452 24834
rect 18396 24770 18452 24782
rect 16492 24658 16548 24668
rect 18508 24500 18564 24510
rect 18508 24406 18564 24444
rect 18620 24052 18676 25454
rect 18844 25506 18900 25518
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18732 24724 18788 24734
rect 18732 24630 18788 24668
rect 15260 23436 15428 23492
rect 18396 23996 18676 24052
rect 15260 23268 15316 23436
rect 15148 22596 15204 22606
rect 15260 22596 15316 23212
rect 17388 23268 17444 23278
rect 17388 23174 17444 23212
rect 17724 23156 17780 23166
rect 17612 23100 17724 23156
rect 15148 22594 15316 22596
rect 15148 22542 15150 22594
rect 15202 22542 15316 22594
rect 15148 22540 15316 22542
rect 15372 23042 15428 23054
rect 15372 22990 15374 23042
rect 15426 22990 15428 23042
rect 15148 22530 15204 22540
rect 15372 22372 15428 22990
rect 16380 22484 16436 22494
rect 16380 22390 16436 22428
rect 15372 22306 15428 22316
rect 16156 22372 16212 22382
rect 16156 22278 16212 22316
rect 17388 22372 17444 22382
rect 17388 22278 17444 22316
rect 15484 22146 15540 22158
rect 15820 22148 15876 22158
rect 15484 22094 15486 22146
rect 15538 22094 15540 22146
rect 15372 21812 15428 21822
rect 15036 21810 15428 21812
rect 15036 21758 15374 21810
rect 15426 21758 15428 21810
rect 15036 21756 15428 21758
rect 14700 21476 14756 21486
rect 14588 21474 14756 21476
rect 14588 21422 14702 21474
rect 14754 21422 14756 21474
rect 14588 21420 14756 21422
rect 14252 21410 14308 21420
rect 14588 20580 14644 20590
rect 14476 20578 14644 20580
rect 14476 20526 14590 20578
rect 14642 20526 14644 20578
rect 14476 20524 14644 20526
rect 14476 20188 14532 20524
rect 14588 20514 14644 20524
rect 11340 19966 11342 20018
rect 11394 19966 11396 20018
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 11340 19012 11396 19966
rect 14140 20132 14532 20188
rect 14140 20020 14196 20132
rect 12012 19908 12068 19918
rect 12012 19814 12068 19852
rect 14140 19906 14196 19964
rect 14588 20130 14644 20142
rect 14588 20078 14590 20130
rect 14642 20078 14644 20130
rect 14140 19854 14142 19906
rect 14194 19854 14196 19906
rect 14140 19842 14196 19854
rect 14476 19908 14532 19918
rect 14476 19814 14532 19852
rect 14588 19460 14644 20078
rect 14588 19394 14644 19404
rect 14476 19234 14532 19246
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 13804 19012 13860 19022
rect 11340 18946 11396 18956
rect 13580 18956 13804 19012
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 10668 18452 10724 18462
rect 10668 18338 10724 18396
rect 13580 18450 13636 18956
rect 13804 18918 13860 18956
rect 14028 18900 14084 18910
rect 14028 18674 14084 18844
rect 14028 18622 14030 18674
rect 14082 18622 14084 18674
rect 14028 18610 14084 18622
rect 13580 18398 13582 18450
rect 13634 18398 13636 18450
rect 10668 18286 10670 18338
rect 10722 18286 10724 18338
rect 10668 18274 10724 18286
rect 12348 18340 12404 18350
rect 12796 18340 12852 18350
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 12348 17778 12404 18284
rect 12460 18338 12852 18340
rect 12460 18286 12798 18338
rect 12850 18286 12852 18338
rect 12460 18284 12852 18286
rect 12460 17890 12516 18284
rect 12796 18274 12852 18284
rect 12460 17838 12462 17890
rect 12514 17838 12516 17890
rect 12460 17826 12516 17838
rect 12348 17726 12350 17778
rect 12402 17726 12404 17778
rect 12348 17714 12404 17726
rect 13580 17666 13636 18398
rect 14252 18562 14308 18574
rect 14252 18510 14254 18562
rect 14306 18510 14308 18562
rect 14252 18452 14308 18510
rect 14252 18386 14308 18396
rect 14476 18564 14532 19182
rect 14588 19122 14644 19134
rect 14588 19070 14590 19122
rect 14642 19070 14644 19122
rect 14588 18900 14644 19070
rect 14700 19012 14756 21420
rect 15036 20188 15092 21756
rect 15372 21746 15428 21756
rect 15148 20916 15204 20926
rect 15148 20822 15204 20860
rect 15484 20692 15540 22094
rect 15484 20626 15540 20636
rect 15708 22146 15876 22148
rect 15708 22094 15822 22146
rect 15874 22094 15876 22146
rect 15708 22092 15876 22094
rect 15708 21810 15764 22092
rect 15820 22082 15876 22092
rect 15708 21758 15710 21810
rect 15762 21758 15764 21810
rect 14924 20132 15092 20188
rect 15708 20188 15764 21758
rect 17612 21810 17668 23100
rect 17724 23062 17780 23100
rect 18172 23154 18228 23166
rect 18172 23102 18174 23154
rect 18226 23102 18228 23154
rect 18172 22484 18228 23102
rect 18172 22418 18228 22428
rect 17836 22258 17892 22270
rect 17836 22206 17838 22258
rect 17890 22206 17892 22258
rect 17836 21924 17892 22206
rect 18396 22148 18452 23996
rect 18508 23826 18564 23838
rect 18508 23774 18510 23826
rect 18562 23774 18564 23826
rect 18508 22372 18564 23774
rect 18620 23716 18676 23726
rect 18844 23716 18900 25454
rect 18956 25508 19012 25518
rect 19292 25508 19348 25564
rect 20188 25618 20468 25620
rect 20188 25566 20190 25618
rect 20242 25566 20468 25618
rect 20188 25564 20468 25566
rect 20524 26404 20580 26414
rect 20188 25554 20244 25564
rect 19852 25508 19908 25518
rect 19292 25506 19908 25508
rect 19292 25454 19854 25506
rect 19906 25454 19908 25506
rect 19292 25452 19908 25454
rect 18956 24948 19012 25452
rect 19852 25442 19908 25452
rect 19180 25394 19236 25406
rect 19180 25342 19182 25394
rect 19234 25342 19236 25394
rect 19180 25284 19236 25342
rect 20076 25396 20132 25406
rect 20076 25302 20132 25340
rect 20188 25394 20244 25406
rect 20188 25342 20190 25394
rect 20242 25342 20244 25394
rect 19236 25228 19348 25284
rect 19180 25218 19236 25228
rect 18956 24722 19012 24892
rect 18956 24670 18958 24722
rect 19010 24670 19012 24722
rect 18956 24658 19012 24670
rect 19180 24724 19236 24734
rect 18620 23714 18900 23716
rect 18620 23662 18622 23714
rect 18674 23662 18900 23714
rect 18620 23660 18900 23662
rect 18956 24500 19012 24510
rect 18956 23714 19012 24444
rect 18956 23662 18958 23714
rect 19010 23662 19012 23714
rect 18620 23650 18676 23660
rect 18620 23268 18676 23278
rect 18620 23042 18676 23212
rect 18620 22990 18622 23042
rect 18674 22990 18676 23042
rect 18620 22596 18676 22990
rect 18732 23044 18788 23660
rect 18956 23268 19012 23662
rect 18956 23202 19012 23212
rect 19180 23266 19236 24668
rect 19292 23826 19348 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19292 23774 19294 23826
rect 19346 23774 19348 23826
rect 19292 23762 19348 23774
rect 19628 24388 19684 24398
rect 19628 23378 19684 24332
rect 20188 24388 20244 25342
rect 20188 24322 20244 24332
rect 20300 25396 20356 25406
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23326 19630 23378
rect 19682 23326 19684 23378
rect 19628 23314 19684 23326
rect 20300 23380 20356 25340
rect 20412 24948 20468 24958
rect 20524 24948 20580 26348
rect 20748 26404 20804 26414
rect 20748 26310 20804 26348
rect 20860 26068 20916 26078
rect 20636 26066 20916 26068
rect 20636 26014 20862 26066
rect 20914 26014 20916 26066
rect 20636 26012 20916 26014
rect 20636 25506 20692 26012
rect 20860 26002 20916 26012
rect 22428 25730 22484 26908
rect 22428 25678 22430 25730
rect 22482 25678 22484 25730
rect 22428 25666 22484 25678
rect 22540 26292 22596 26302
rect 20636 25454 20638 25506
rect 20690 25454 20692 25506
rect 20636 25442 20692 25454
rect 22316 25620 22372 25630
rect 22316 25284 22372 25564
rect 22428 25396 22484 25406
rect 22428 25302 22484 25340
rect 22540 25394 22596 26236
rect 22540 25342 22542 25394
rect 22594 25342 22596 25394
rect 22316 25218 22372 25228
rect 22540 25284 22596 25342
rect 22540 25218 22596 25228
rect 22652 25956 22708 25966
rect 20412 24946 20524 24948
rect 20412 24894 20414 24946
rect 20466 24894 20524 24946
rect 20412 24892 20524 24894
rect 20412 24882 20468 24892
rect 20524 24882 20580 24892
rect 21868 24892 22484 24948
rect 20748 24724 20804 24734
rect 20748 24630 20804 24668
rect 20300 23314 20356 23324
rect 20860 23380 20916 23390
rect 20860 23286 20916 23324
rect 19180 23214 19182 23266
rect 19234 23214 19236 23266
rect 19068 23156 19124 23166
rect 19068 23062 19124 23100
rect 18732 22978 18788 22988
rect 19180 22820 19236 23214
rect 19964 23266 20020 23278
rect 19964 23214 19966 23266
rect 20018 23214 20020 23266
rect 19964 23156 20020 23214
rect 19964 23090 20020 23100
rect 20636 23156 20692 23166
rect 18620 22530 18676 22540
rect 18732 22764 19236 22820
rect 19628 23044 19684 23054
rect 18508 22306 18564 22316
rect 18396 22092 18564 22148
rect 17836 21858 17892 21868
rect 18284 21924 18340 21934
rect 17612 21758 17614 21810
rect 17666 21758 17668 21810
rect 17612 21746 17668 21758
rect 17500 21700 17556 21710
rect 17500 21606 17556 21644
rect 17948 21700 18004 21710
rect 17836 21586 17892 21598
rect 17836 21534 17838 21586
rect 17890 21534 17892 21586
rect 16828 21476 16884 21486
rect 16828 21382 16884 21420
rect 17500 20690 17556 20702
rect 17500 20638 17502 20690
rect 17554 20638 17556 20690
rect 14812 19794 14868 19806
rect 14812 19742 14814 19794
rect 14866 19742 14868 19794
rect 14812 19346 14868 19742
rect 14812 19294 14814 19346
rect 14866 19294 14868 19346
rect 14812 19282 14868 19294
rect 14700 18946 14756 18956
rect 14924 19122 14980 20132
rect 15596 20130 15652 20142
rect 15708 20132 16324 20188
rect 15596 20078 15598 20130
rect 15650 20078 15652 20130
rect 15260 20020 15316 20030
rect 15260 19926 15316 19964
rect 15596 19684 15652 20078
rect 16268 20018 16324 20132
rect 16268 19966 16270 20018
rect 16322 19966 16324 20018
rect 16268 19954 16324 19966
rect 16492 19906 16548 19918
rect 16492 19854 16494 19906
rect 16546 19854 16548 19906
rect 15596 19618 15652 19628
rect 15932 19794 15988 19806
rect 15932 19742 15934 19794
rect 15986 19742 15988 19794
rect 15932 19460 15988 19742
rect 15932 19394 15988 19404
rect 16044 19684 16100 19694
rect 16044 19234 16100 19628
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 16044 19170 16100 19182
rect 14924 19070 14926 19122
rect 14978 19070 14980 19122
rect 14588 18834 14644 18844
rect 14700 18788 14756 18798
rect 14476 18450 14532 18508
rect 14588 18564 14644 18574
rect 14700 18564 14756 18732
rect 14588 18562 14756 18564
rect 14588 18510 14590 18562
rect 14642 18510 14756 18562
rect 14588 18508 14756 18510
rect 14588 18498 14644 18508
rect 14476 18398 14478 18450
rect 14530 18398 14532 18450
rect 14476 18386 14532 18398
rect 14140 18340 14196 18350
rect 14140 18246 14196 18284
rect 13580 17614 13582 17666
rect 13634 17614 13636 17666
rect 13580 17602 13636 17614
rect 14252 17554 14308 17566
rect 14252 17502 14254 17554
rect 14306 17502 14308 17554
rect 14252 16996 14308 17502
rect 14252 16930 14308 16940
rect 4284 16884 4340 16894
rect 4284 16790 4340 16828
rect 12460 16884 12516 16894
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16146 1988 16156
rect 12460 15988 12516 16828
rect 14924 16882 14980 19070
rect 16492 19124 16548 19854
rect 17388 19906 17444 19918
rect 17388 19854 17390 19906
rect 17442 19854 17444 19906
rect 16492 19058 16548 19068
rect 17052 19124 17108 19134
rect 15372 19012 15428 19022
rect 15372 18918 15428 18956
rect 15708 19010 15764 19022
rect 15708 18958 15710 19010
rect 15762 18958 15764 19010
rect 15260 18676 15316 18686
rect 15036 16996 15092 17006
rect 15036 16902 15092 16940
rect 15260 16994 15316 18620
rect 15260 16942 15262 16994
rect 15314 16942 15316 16994
rect 15260 16930 15316 16942
rect 15708 18564 15764 18958
rect 16716 19010 16772 19022
rect 16716 18958 16718 19010
rect 16770 18958 16772 19010
rect 16716 18676 16772 18958
rect 16716 18610 16772 18620
rect 16940 19010 16996 19022
rect 16940 18958 16942 19010
rect 16994 18958 16996 19010
rect 14924 16830 14926 16882
rect 14978 16830 14980 16882
rect 14924 16660 14980 16830
rect 14924 16594 14980 16604
rect 15372 16884 15428 16894
rect 12460 15202 12516 15932
rect 15372 15986 15428 16828
rect 15484 16882 15540 16894
rect 15484 16830 15486 16882
rect 15538 16830 15540 16882
rect 15484 16772 15540 16830
rect 15708 16884 15764 18508
rect 16492 18338 16548 18350
rect 16492 18286 16494 18338
rect 16546 18286 16548 18338
rect 16380 17780 16436 17790
rect 16492 17780 16548 18286
rect 16828 18340 16884 18350
rect 16828 18246 16884 18284
rect 16380 17778 16548 17780
rect 16380 17726 16382 17778
rect 16434 17726 16548 17778
rect 16380 17724 16548 17726
rect 16380 17668 16436 17724
rect 16940 17668 16996 18958
rect 17052 17890 17108 19068
rect 17388 19124 17444 19854
rect 17388 19058 17444 19068
rect 17052 17838 17054 17890
rect 17106 17838 17108 17890
rect 17052 17826 17108 17838
rect 17500 19012 17556 20638
rect 17836 20356 17892 21534
rect 17836 20290 17892 20300
rect 17948 20916 18004 21644
rect 18284 21586 18340 21868
rect 18284 21534 18286 21586
rect 18338 21534 18340 21586
rect 18284 21522 18340 21534
rect 17948 20242 18004 20860
rect 17948 20190 17950 20242
rect 18002 20190 18004 20242
rect 17948 20188 18004 20190
rect 17948 20132 18116 20188
rect 17948 19458 18004 19470
rect 17948 19406 17950 19458
rect 18002 19406 18004 19458
rect 17612 19234 17668 19246
rect 17612 19182 17614 19234
rect 17666 19182 17668 19234
rect 17612 19124 17668 19182
rect 17612 19058 17668 19068
rect 17948 19124 18004 19406
rect 17500 18338 17556 18956
rect 17836 19012 17892 19022
rect 17500 18286 17502 18338
rect 17554 18286 17556 18338
rect 17388 17668 17444 17678
rect 16940 17666 17444 17668
rect 16940 17614 17390 17666
rect 17442 17614 17444 17666
rect 16940 17612 17444 17614
rect 16380 17602 16436 17612
rect 15708 16818 15764 16828
rect 16828 17444 16884 17454
rect 16828 16882 16884 17388
rect 17164 17442 17220 17454
rect 17164 17390 17166 17442
rect 17218 17390 17220 17442
rect 17164 16996 17220 17390
rect 17388 17108 17444 17612
rect 17500 17220 17556 18286
rect 17724 18788 17780 18798
rect 17724 18340 17780 18732
rect 17836 18674 17892 18956
rect 17948 18788 18004 19068
rect 17948 18722 18004 18732
rect 17836 18622 17838 18674
rect 17890 18622 17892 18674
rect 17836 18610 17892 18622
rect 17948 18452 18004 18462
rect 17724 18284 17892 18340
rect 17724 17668 17780 17678
rect 17724 17574 17780 17612
rect 17500 17164 17780 17220
rect 17388 17052 17668 17108
rect 17164 16930 17220 16940
rect 16828 16830 16830 16882
rect 16882 16830 16884 16882
rect 16828 16818 16884 16830
rect 17388 16884 17444 16894
rect 17388 16790 17444 16828
rect 17612 16882 17668 17052
rect 17612 16830 17614 16882
rect 17666 16830 17668 16882
rect 15484 16706 15540 16716
rect 16268 16772 16324 16782
rect 15820 16548 15876 16558
rect 15820 16098 15876 16492
rect 15820 16046 15822 16098
rect 15874 16046 15876 16098
rect 15820 16034 15876 16046
rect 15372 15934 15374 15986
rect 15426 15934 15428 15986
rect 15372 15922 15428 15934
rect 15596 15988 15652 15998
rect 15596 15894 15652 15932
rect 15708 15874 15764 15886
rect 15708 15822 15710 15874
rect 15762 15822 15764 15874
rect 15708 15428 15764 15822
rect 15708 15372 16100 15428
rect 15372 15314 15428 15326
rect 15372 15262 15374 15314
rect 15426 15262 15428 15314
rect 12460 15150 12462 15202
rect 12514 15150 12516 15202
rect 12460 15138 12516 15150
rect 14028 15204 14084 15214
rect 14588 15204 14644 15214
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14028 14642 14084 15148
rect 14140 15202 14644 15204
rect 14140 15150 14590 15202
rect 14642 15150 14644 15202
rect 14140 15148 14644 15150
rect 14140 14754 14196 15148
rect 14588 15138 14644 15148
rect 14140 14702 14142 14754
rect 14194 14702 14196 14754
rect 14140 14690 14196 14702
rect 14028 14590 14030 14642
rect 14082 14590 14084 14642
rect 14028 14578 14084 14590
rect 15372 14308 15428 15262
rect 16044 15314 16100 15372
rect 16268 15426 16324 16716
rect 16604 16772 16660 16782
rect 16604 16678 16660 16716
rect 17276 16772 17332 16782
rect 16492 16660 16548 16670
rect 16492 16566 16548 16604
rect 17276 16098 17332 16716
rect 17500 16770 17556 16782
rect 17500 16718 17502 16770
rect 17554 16718 17556 16770
rect 17500 16324 17556 16718
rect 17612 16548 17668 16830
rect 17724 16884 17780 17164
rect 17836 17106 17892 18284
rect 17948 17556 18004 18396
rect 18060 17892 18116 20132
rect 18172 19122 18228 19134
rect 18172 19070 18174 19122
rect 18226 19070 18228 19122
rect 18172 18450 18228 19070
rect 18508 18676 18564 22092
rect 18732 21586 18788 22764
rect 18956 22484 19012 22494
rect 18956 22390 19012 22428
rect 19516 22484 19572 22494
rect 19068 22372 19124 22382
rect 19068 21588 19124 22316
rect 18732 21534 18734 21586
rect 18786 21534 18788 21586
rect 18732 20244 18788 21534
rect 18956 21532 19124 21588
rect 19180 22370 19236 22382
rect 19180 22318 19182 22370
rect 19234 22318 19236 22370
rect 19180 21924 19236 22318
rect 19292 22372 19348 22382
rect 19292 22146 19348 22316
rect 19292 22094 19294 22146
rect 19346 22094 19348 22146
rect 19292 22082 19348 22094
rect 18956 20188 19012 21532
rect 18732 20178 18788 20188
rect 18844 20132 19012 20188
rect 19068 20244 19124 20254
rect 18620 20018 18676 20030
rect 18620 19966 18622 20018
rect 18674 19966 18676 20018
rect 18620 19684 18676 19966
rect 18620 19618 18676 19628
rect 18732 19796 18788 19806
rect 18508 18610 18564 18620
rect 18172 18398 18174 18450
rect 18226 18398 18228 18450
rect 18172 18340 18228 18398
rect 18620 18452 18676 18462
rect 18620 18358 18676 18396
rect 18172 18274 18228 18284
rect 18508 18340 18564 18350
rect 18060 17826 18116 17836
rect 18060 17556 18116 17566
rect 17948 17554 18116 17556
rect 17948 17502 18062 17554
rect 18114 17502 18116 17554
rect 17948 17500 18116 17502
rect 18060 17490 18116 17500
rect 18396 17444 18452 17454
rect 18396 17350 18452 17388
rect 17836 17054 17838 17106
rect 17890 17054 17892 17106
rect 17836 17042 17892 17054
rect 18284 16994 18340 17006
rect 18284 16942 18286 16994
rect 18338 16942 18340 16994
rect 18060 16884 18116 16894
rect 17724 16828 18004 16884
rect 17612 16482 17668 16492
rect 17836 16324 17892 16334
rect 17500 16322 17892 16324
rect 17500 16270 17838 16322
rect 17890 16270 17892 16322
rect 17500 16268 17892 16270
rect 17836 16258 17892 16268
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 17276 16034 17332 16046
rect 16268 15374 16270 15426
rect 16322 15374 16324 15426
rect 16268 15362 16324 15374
rect 17612 15986 17668 15998
rect 17612 15934 17614 15986
rect 17666 15934 17668 15986
rect 16044 15262 16046 15314
rect 16098 15262 16100 15314
rect 16044 15250 16100 15262
rect 15708 15204 15764 15214
rect 15708 15110 15764 15148
rect 17612 15204 17668 15934
rect 17612 15138 17668 15148
rect 17836 14532 17892 14542
rect 17948 14532 18004 16828
rect 18060 16210 18116 16828
rect 18284 16548 18340 16942
rect 18508 16882 18564 18284
rect 18732 17780 18788 19740
rect 18508 16830 18510 16882
rect 18562 16830 18564 16882
rect 18508 16818 18564 16830
rect 18620 17724 18788 17780
rect 18284 16482 18340 16492
rect 18060 16158 18062 16210
rect 18114 16158 18116 16210
rect 18060 16146 18116 16158
rect 18284 15988 18340 15998
rect 18284 15986 18564 15988
rect 18284 15934 18286 15986
rect 18338 15934 18564 15986
rect 18284 15932 18564 15934
rect 18284 15922 18340 15932
rect 17836 14530 18004 14532
rect 17836 14478 17838 14530
rect 17890 14478 18004 14530
rect 17836 14476 18004 14478
rect 18172 15874 18228 15886
rect 18172 15822 18174 15874
rect 18226 15822 18228 15874
rect 15596 14308 15652 14318
rect 15372 14252 15596 14308
rect 15596 14214 15652 14252
rect 17500 14308 17556 14318
rect 17836 14308 17892 14476
rect 17556 14252 17892 14308
rect 17500 13748 17556 14252
rect 18172 13858 18228 15822
rect 18508 15538 18564 15932
rect 18508 15486 18510 15538
rect 18562 15486 18564 15538
rect 18508 15474 18564 15486
rect 18620 15540 18676 17724
rect 18732 17442 18788 17454
rect 18732 17390 18734 17442
rect 18786 17390 18788 17442
rect 18732 17220 18788 17390
rect 18844 17444 18900 20132
rect 19068 19234 19124 20188
rect 19180 20020 19236 21868
rect 19404 21586 19460 21598
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 21476 19460 21534
rect 19404 21410 19460 21420
rect 19404 20356 19460 20366
rect 19180 19954 19236 19964
rect 19292 20018 19348 20030
rect 19292 19966 19294 20018
rect 19346 19966 19348 20018
rect 19068 19182 19070 19234
rect 19122 19182 19124 19234
rect 19068 19170 19124 19182
rect 19292 18564 19348 19966
rect 19180 18508 19348 18564
rect 18956 18340 19012 18350
rect 19180 18340 19236 18508
rect 19404 18452 19460 20300
rect 19516 19234 19572 22428
rect 19516 19182 19518 19234
rect 19570 19182 19572 19234
rect 19516 19170 19572 19182
rect 19404 18358 19460 18396
rect 18956 18338 19236 18340
rect 18956 18286 18958 18338
rect 19010 18286 19236 18338
rect 18956 18284 19236 18286
rect 19292 18340 19348 18350
rect 18956 17668 19012 18284
rect 18956 17602 19012 17612
rect 19068 17892 19124 17902
rect 19068 17666 19124 17836
rect 19292 17890 19348 18284
rect 19292 17838 19294 17890
rect 19346 17838 19348 17890
rect 19292 17826 19348 17838
rect 19516 17892 19572 17902
rect 19628 17892 19684 22988
rect 20188 22258 20244 22270
rect 20188 22206 20190 22258
rect 20242 22206 20244 22258
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 22206
rect 20636 22260 20692 23100
rect 21868 23154 21924 24892
rect 21868 23102 21870 23154
rect 21922 23102 21924 23154
rect 21868 23090 21924 23102
rect 22316 24724 22372 24734
rect 22428 24724 22484 24892
rect 22652 24946 22708 25900
rect 22876 25508 22932 27020
rect 22988 27010 23044 27020
rect 23660 26964 23716 27806
rect 23772 27634 23828 27646
rect 23772 27582 23774 27634
rect 23826 27582 23828 27634
rect 23772 27186 23828 27582
rect 23772 27134 23774 27186
rect 23826 27134 23828 27186
rect 23772 27122 23828 27134
rect 23660 26898 23716 26908
rect 23884 26516 23940 26526
rect 23884 26422 23940 26460
rect 23436 26292 23492 26302
rect 23324 26290 23492 26292
rect 23324 26238 23438 26290
rect 23490 26238 23492 26290
rect 23324 26236 23492 26238
rect 22988 26180 23044 26190
rect 22988 26086 23044 26124
rect 23100 26068 23156 26078
rect 23100 25974 23156 26012
rect 22652 24894 22654 24946
rect 22706 24894 22708 24946
rect 22652 24882 22708 24894
rect 22764 25506 22932 25508
rect 22764 25454 22878 25506
rect 22930 25454 22932 25506
rect 22764 25452 22932 25454
rect 22764 24724 22820 25452
rect 22876 25442 22932 25452
rect 23324 25620 23380 26236
rect 23436 26226 23492 26236
rect 23660 26292 23716 26302
rect 23660 26198 23716 26236
rect 23996 26292 24052 26302
rect 23772 26180 23828 26190
rect 23772 26086 23828 26124
rect 22428 24668 22820 24724
rect 21308 22484 21364 22494
rect 21308 22390 21364 22428
rect 22316 22372 22372 24668
rect 22652 23826 22708 23838
rect 22652 23774 22654 23826
rect 22706 23774 22708 23826
rect 22540 23714 22596 23726
rect 22540 23662 22542 23714
rect 22594 23662 22596 23714
rect 22540 23042 22596 23662
rect 22652 23492 22708 23774
rect 22652 23426 22708 23436
rect 22540 22990 22542 23042
rect 22594 22990 22596 23042
rect 22540 22978 22596 22990
rect 21980 22370 22372 22372
rect 21980 22318 22318 22370
rect 22370 22318 22372 22370
rect 21980 22316 22372 22318
rect 20636 22194 20692 22204
rect 21644 22260 21700 22270
rect 21700 22204 21924 22260
rect 21644 22166 21700 22204
rect 20076 21756 20244 21812
rect 20076 21700 20132 21756
rect 20076 21634 20132 21644
rect 20076 21476 20132 21486
rect 20076 20802 20132 21420
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 21420 20802 21476 20814
rect 21420 20750 21422 20802
rect 21474 20750 21476 20802
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 21420 20244 21476 20750
rect 21644 20802 21700 20814
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21420 20178 21476 20188
rect 21532 20692 21588 20702
rect 19852 20130 19908 20142
rect 19852 20078 19854 20130
rect 19906 20078 19908 20130
rect 19740 19796 19796 19806
rect 19852 19796 19908 20078
rect 19796 19740 19908 19796
rect 20412 20020 20468 20030
rect 19740 19730 19796 19740
rect 20300 19684 20356 19694
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20300 18338 20356 19628
rect 20412 18450 20468 19964
rect 21308 20020 21364 20030
rect 21308 19926 21364 19964
rect 21532 19458 21588 20636
rect 21644 19684 21700 20750
rect 21868 20130 21924 22204
rect 21980 21026 22036 22316
rect 22316 22306 22372 22316
rect 22652 22260 22708 22270
rect 22652 22166 22708 22204
rect 21980 20974 21982 21026
rect 22034 20974 22036 21026
rect 21980 20962 22036 20974
rect 22652 21028 22708 21038
rect 22652 20934 22708 20972
rect 22764 20916 22820 24668
rect 22988 22260 23044 22270
rect 22988 22258 23156 22260
rect 22988 22206 22990 22258
rect 23042 22206 23156 22258
rect 22988 22204 23156 22206
rect 22988 22194 23044 22204
rect 22652 20804 22708 20814
rect 22316 20692 22372 20702
rect 22316 20598 22372 20636
rect 22540 20244 22596 20254
rect 22652 20244 22708 20748
rect 22540 20242 22708 20244
rect 22540 20190 22542 20242
rect 22594 20190 22708 20242
rect 22540 20188 22708 20190
rect 22764 20188 22820 20860
rect 21868 20078 21870 20130
rect 21922 20078 21924 20130
rect 21868 20066 21924 20078
rect 22204 20132 22596 20188
rect 22764 20132 22932 20188
rect 21644 19618 21700 19628
rect 21532 19406 21534 19458
rect 21586 19406 21588 19458
rect 21532 19394 21588 19406
rect 21756 19460 21812 19470
rect 21756 19366 21812 19404
rect 22092 19346 22148 19358
rect 22092 19294 22094 19346
rect 22146 19294 22148 19346
rect 22092 18788 22148 19294
rect 22204 19234 22260 20132
rect 22204 19182 22206 19234
rect 22258 19182 22260 19234
rect 22204 19170 22260 19182
rect 22876 19234 22932 20132
rect 22876 19182 22878 19234
rect 22930 19182 22932 19234
rect 22316 19122 22372 19134
rect 22316 19070 22318 19122
rect 22370 19070 22372 19122
rect 22316 19012 22372 19070
rect 22316 18946 22372 18956
rect 22092 18732 22708 18788
rect 20412 18398 20414 18450
rect 20466 18398 20468 18450
rect 20412 18386 20468 18398
rect 20860 18452 20916 18462
rect 20300 18286 20302 18338
rect 20354 18286 20356 18338
rect 20300 18274 20356 18286
rect 19516 17890 19628 17892
rect 19516 17838 19518 17890
rect 19570 17838 19628 17890
rect 19516 17836 19628 17838
rect 19516 17826 19572 17836
rect 19628 17798 19684 17836
rect 20412 18226 20468 18238
rect 20412 18174 20414 18226
rect 20466 18174 20468 18226
rect 19068 17614 19070 17666
rect 19122 17614 19124 17666
rect 19068 17602 19124 17614
rect 19628 17556 19684 17566
rect 19628 17462 19684 17500
rect 18844 17388 19572 17444
rect 18732 16884 18788 17164
rect 18732 16818 18788 16828
rect 19516 16772 19572 17388
rect 19628 17332 19684 17342
rect 19628 17108 19684 17276
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 19628 17106 19908 17108
rect 19628 17054 19854 17106
rect 19906 17054 19908 17106
rect 19628 17052 19908 17054
rect 19852 17042 19908 17052
rect 19740 16884 19796 16894
rect 19628 16772 19684 16782
rect 19516 16770 19684 16772
rect 19516 16718 19630 16770
rect 19682 16718 19684 16770
rect 19516 16716 19684 16718
rect 19628 16706 19684 16716
rect 19740 15988 19796 16828
rect 19964 16660 20020 16670
rect 20076 16660 20132 16670
rect 19964 16658 20076 16660
rect 19964 16606 19966 16658
rect 20018 16606 20076 16658
rect 19964 16604 20076 16606
rect 20132 16604 20244 16660
rect 19964 16594 20020 16604
rect 20076 16566 20132 16604
rect 19628 15932 19796 15988
rect 18732 15540 18788 15550
rect 18620 15484 18732 15540
rect 18732 15474 18788 15484
rect 19292 15428 19348 15438
rect 19292 15426 19572 15428
rect 19292 15374 19294 15426
rect 19346 15374 19572 15426
rect 19292 15372 19572 15374
rect 19292 15362 19348 15372
rect 18620 15316 18676 15326
rect 18956 15316 19012 15326
rect 18172 13806 18174 13858
rect 18226 13806 18228 13858
rect 18172 13794 18228 13806
rect 18508 15314 19012 15316
rect 18508 15262 18622 15314
rect 18674 15262 18958 15314
rect 19010 15262 19012 15314
rect 18508 15260 19012 15262
rect 17500 13654 17556 13692
rect 18508 13524 18564 15260
rect 18620 15250 18676 15260
rect 18956 15250 19012 15260
rect 18732 14644 18788 14654
rect 18620 14588 18732 14644
rect 18620 14530 18676 14588
rect 18732 14578 18788 14588
rect 18620 14478 18622 14530
rect 18674 14478 18676 14530
rect 18620 14466 18676 14478
rect 18508 13458 18564 13468
rect 19404 13524 19460 13534
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 18844 3666 18900 3678
rect 18844 3614 18846 3666
rect 18898 3614 18900 3666
rect 18844 800 18900 3614
rect 19404 3556 19460 13468
rect 19516 8428 19572 15372
rect 19628 15316 19684 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15540 20244 16604
rect 20412 16212 20468 18174
rect 20860 17556 20916 18396
rect 22316 18450 22372 18462
rect 22316 18398 22318 18450
rect 22370 18398 22372 18450
rect 22204 17892 22260 17902
rect 21756 17668 21812 17678
rect 21868 17668 21924 17678
rect 21756 17666 21868 17668
rect 21756 17614 21758 17666
rect 21810 17614 21868 17666
rect 21756 17612 21868 17614
rect 21756 17602 21812 17612
rect 20860 16994 20916 17500
rect 21420 17108 21476 17118
rect 21420 17014 21476 17052
rect 20860 16942 20862 16994
rect 20914 16942 20916 16994
rect 20860 16930 20916 16942
rect 21084 16660 21140 16670
rect 21084 16566 21140 16604
rect 20412 16146 20468 16156
rect 19964 15484 20244 15540
rect 19740 15316 19796 15326
rect 19628 15314 19796 15316
rect 19628 15262 19742 15314
rect 19794 15262 19796 15314
rect 19628 15260 19796 15262
rect 19740 15250 19796 15260
rect 19964 15314 20020 15484
rect 20636 15428 20692 15438
rect 20412 15426 20692 15428
rect 20412 15374 20638 15426
rect 20690 15374 20692 15426
rect 20412 15372 20692 15374
rect 19964 15262 19966 15314
rect 20018 15262 20020 15314
rect 19964 15250 20020 15262
rect 20188 15316 20244 15326
rect 20412 15316 20468 15372
rect 20636 15362 20692 15372
rect 20748 15426 20804 15438
rect 20748 15374 20750 15426
rect 20802 15374 20804 15426
rect 20188 15314 20468 15316
rect 20188 15262 20190 15314
rect 20242 15262 20468 15314
rect 20188 15260 20468 15262
rect 20188 15250 20244 15260
rect 20524 15204 20580 15214
rect 20524 15110 20580 15148
rect 19628 15090 19684 15102
rect 19628 15038 19630 15090
rect 19682 15038 19684 15090
rect 19628 14644 19684 15038
rect 20748 14644 20804 15374
rect 21868 15314 21924 17612
rect 22204 16994 22260 17836
rect 22316 17108 22372 18398
rect 22652 18450 22708 18732
rect 22652 18398 22654 18450
rect 22706 18398 22708 18450
rect 22652 18386 22708 18398
rect 22540 18338 22596 18350
rect 22540 18286 22542 18338
rect 22594 18286 22596 18338
rect 22428 17780 22484 17790
rect 22540 17780 22596 18286
rect 22428 17778 22596 17780
rect 22428 17726 22430 17778
rect 22482 17726 22596 17778
rect 22428 17724 22596 17726
rect 22428 17714 22484 17724
rect 22876 17668 22932 19182
rect 22876 17602 22932 17612
rect 22988 20132 23044 20142
rect 22988 18450 23044 20076
rect 23100 19012 23156 22204
rect 23212 22258 23268 22270
rect 23212 22206 23214 22258
rect 23266 22206 23268 22258
rect 23212 21028 23268 22206
rect 23324 21700 23380 25564
rect 23660 26068 23716 26078
rect 23660 25618 23716 26012
rect 23996 25956 24052 26236
rect 24332 26068 24388 27916
rect 24556 27188 24612 27198
rect 24556 26514 24612 27132
rect 24556 26462 24558 26514
rect 24610 26462 24612 26514
rect 24556 26450 24612 26462
rect 25788 26516 25844 31892
rect 25900 27188 25956 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25900 27094 25956 27132
rect 24444 26292 24500 26302
rect 24444 26198 24500 26236
rect 24556 26068 24612 26078
rect 24332 26066 24612 26068
rect 24332 26014 24558 26066
rect 24610 26014 24612 26066
rect 24332 26012 24612 26014
rect 24556 26002 24612 26012
rect 23996 25890 24052 25900
rect 23660 25566 23662 25618
rect 23714 25566 23716 25618
rect 23660 25554 23716 25566
rect 25788 25618 25844 26460
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 25788 25566 25790 25618
rect 25842 25566 25844 25618
rect 25788 25554 25844 25566
rect 23436 25284 23492 25294
rect 23436 22370 23492 25228
rect 26572 24722 26628 24734
rect 26572 24670 26574 24722
rect 26626 24670 26628 24722
rect 25900 24388 25956 24398
rect 25900 23716 25956 24332
rect 24556 23492 24612 23502
rect 24444 22932 24500 22942
rect 23436 22318 23438 22370
rect 23490 22318 23492 22370
rect 23436 21812 23492 22318
rect 23660 22428 24052 22484
rect 23660 22370 23716 22428
rect 23660 22318 23662 22370
rect 23714 22318 23716 22370
rect 23660 22306 23716 22318
rect 23884 22258 23940 22270
rect 23884 22206 23886 22258
rect 23938 22206 23940 22258
rect 23772 22148 23828 22158
rect 23660 22146 23828 22148
rect 23660 22094 23774 22146
rect 23826 22094 23828 22146
rect 23660 22092 23828 22094
rect 23436 21756 23604 21812
rect 23324 21644 23492 21700
rect 23212 20962 23268 20972
rect 23324 21476 23380 21486
rect 23324 20802 23380 21420
rect 23324 20750 23326 20802
rect 23378 20750 23380 20802
rect 23324 20738 23380 20750
rect 23436 20188 23492 21644
rect 23100 18946 23156 18956
rect 23324 20132 23492 20188
rect 23324 18676 23380 20132
rect 23548 20018 23604 21756
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 23548 18676 23604 19966
rect 23660 19346 23716 22092
rect 23772 22082 23828 22092
rect 23884 21252 23940 22206
rect 23884 21186 23940 21196
rect 23996 20188 24052 22428
rect 24444 22370 24500 22876
rect 24444 22318 24446 22370
rect 24498 22318 24500 22370
rect 24444 22306 24500 22318
rect 24220 22258 24276 22270
rect 24220 22206 24222 22258
rect 24274 22206 24276 22258
rect 24220 20804 24276 22206
rect 24556 22146 24612 23436
rect 24668 23042 24724 23054
rect 24668 22990 24670 23042
rect 24722 22990 24724 23042
rect 24668 22932 24724 22990
rect 24668 22866 24724 22876
rect 24780 22260 24836 22270
rect 24780 22166 24836 22204
rect 24556 22094 24558 22146
rect 24610 22094 24612 22146
rect 24556 22082 24612 22094
rect 24220 20738 24276 20748
rect 25228 21252 25284 21262
rect 23772 20132 23828 20142
rect 23996 20132 24500 20188
rect 23772 20038 23828 20076
rect 23660 19294 23662 19346
rect 23714 19294 23716 19346
rect 23660 19282 23716 19294
rect 23660 18676 23716 18686
rect 23324 18620 23492 18676
rect 23548 18674 23716 18676
rect 23548 18622 23662 18674
rect 23714 18622 23716 18674
rect 23548 18620 23716 18622
rect 22988 18398 22990 18450
rect 23042 18398 23044 18450
rect 22652 17220 22708 17230
rect 22540 17108 22596 17118
rect 22316 17106 22596 17108
rect 22316 17054 22542 17106
rect 22594 17054 22596 17106
rect 22316 17052 22596 17054
rect 22540 17042 22596 17052
rect 22652 17106 22708 17164
rect 22652 17054 22654 17106
rect 22706 17054 22708 17106
rect 22652 17042 22708 17054
rect 22204 16942 22206 16994
rect 22258 16942 22260 16994
rect 22204 16930 22260 16942
rect 22764 16996 22820 17006
rect 22764 16902 22820 16940
rect 22428 16884 22484 16894
rect 22428 16790 22484 16828
rect 22988 16660 23044 18398
rect 23324 18452 23380 18462
rect 23324 18358 23380 18396
rect 23436 17106 23492 18620
rect 23660 18610 23716 18620
rect 23436 17054 23438 17106
rect 23490 17054 23492 17106
rect 23436 17042 23492 17054
rect 23660 17108 23716 17118
rect 24220 17108 24276 17118
rect 23660 17106 24276 17108
rect 23660 17054 23662 17106
rect 23714 17054 24222 17106
rect 24274 17054 24276 17106
rect 23660 17052 24276 17054
rect 23660 17042 23716 17052
rect 23212 16884 23268 16894
rect 23212 16790 23268 16828
rect 23548 16770 23604 16782
rect 23548 16718 23550 16770
rect 23602 16718 23604 16770
rect 23548 16660 23604 16718
rect 22988 16604 23268 16660
rect 23100 16212 23156 16222
rect 22540 16210 23156 16212
rect 22540 16158 23102 16210
rect 23154 16158 23156 16210
rect 22540 16156 23156 16158
rect 22540 15426 22596 16156
rect 23100 16146 23156 16156
rect 23212 15986 23268 16604
rect 23436 16604 23604 16660
rect 23436 16322 23492 16604
rect 23436 16270 23438 16322
rect 23490 16270 23492 16322
rect 23436 16258 23492 16270
rect 23772 16322 23828 17052
rect 24220 17042 24276 17052
rect 24444 16996 24500 20132
rect 25228 20130 25284 21196
rect 25340 20916 25396 20926
rect 25340 20822 25396 20860
rect 25228 20078 25230 20130
rect 25282 20078 25284 20130
rect 25228 20066 25284 20078
rect 25340 19906 25396 19918
rect 25340 19854 25342 19906
rect 25394 19854 25396 19906
rect 25340 19348 25396 19854
rect 25788 19348 25844 19358
rect 25340 19292 25788 19348
rect 25788 19254 25844 19292
rect 25900 19236 25956 23660
rect 26572 21588 26628 24670
rect 28252 24724 28308 24734
rect 27356 24610 27412 24622
rect 27356 24558 27358 24610
rect 27410 24558 27412 24610
rect 27356 24164 27412 24558
rect 27468 24164 27524 24174
rect 27356 24162 27524 24164
rect 27356 24110 27470 24162
rect 27522 24110 27524 24162
rect 27356 24108 27524 24110
rect 27468 24098 27524 24108
rect 27580 23828 27636 23838
rect 28028 23828 28084 23838
rect 27580 23826 28084 23828
rect 27580 23774 27582 23826
rect 27634 23774 28030 23826
rect 28082 23774 28084 23826
rect 27580 23772 28084 23774
rect 27580 23762 27636 23772
rect 28028 23762 28084 23772
rect 28252 23826 28308 24668
rect 29484 24724 29540 24734
rect 29484 24610 29540 24668
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 29484 24558 29486 24610
rect 29538 24558 29540 24610
rect 29484 24546 29540 24558
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23938 37716 23950
rect 37660 23886 37662 23938
rect 37714 23886 37716 23938
rect 28252 23774 28254 23826
rect 28306 23774 28308 23826
rect 28252 23762 28308 23774
rect 28364 23826 28420 23838
rect 28364 23774 28366 23826
rect 28418 23774 28420 23826
rect 27468 23716 27524 23726
rect 27468 23622 27524 23660
rect 27356 23268 27412 23278
rect 27132 23154 27188 23166
rect 27132 23102 27134 23154
rect 27186 23102 27188 23154
rect 26572 20916 26628 21532
rect 26572 20850 26628 20860
rect 27020 22484 27076 22494
rect 26684 19236 26740 19246
rect 25900 19234 26740 19236
rect 25900 19182 26686 19234
rect 26738 19182 26740 19234
rect 25900 19180 26740 19182
rect 25900 18562 25956 19180
rect 26684 19170 26740 19180
rect 26124 19012 26180 19022
rect 26124 18674 26180 18956
rect 26908 19012 26964 19022
rect 26908 18918 26964 18956
rect 26124 18622 26126 18674
rect 26178 18622 26180 18674
rect 26124 18610 26180 18622
rect 26348 18788 26404 18798
rect 25900 18510 25902 18562
rect 25954 18510 25956 18562
rect 25900 18498 25956 18510
rect 26348 18562 26404 18732
rect 26348 18510 26350 18562
rect 26402 18510 26404 18562
rect 25676 18004 25732 18014
rect 24556 17778 24612 17790
rect 24556 17726 24558 17778
rect 24610 17726 24612 17778
rect 24556 17220 24612 17726
rect 24612 17164 24836 17220
rect 24556 17154 24612 17164
rect 24556 16996 24612 17006
rect 24444 16994 24612 16996
rect 24444 16942 24558 16994
rect 24610 16942 24612 16994
rect 24444 16940 24612 16942
rect 23884 16884 23940 16894
rect 24556 16884 24612 16940
rect 23884 16882 24052 16884
rect 23884 16830 23886 16882
rect 23938 16830 24052 16882
rect 23884 16828 24052 16830
rect 23884 16818 23940 16828
rect 23772 16270 23774 16322
rect 23826 16270 23828 16322
rect 23772 16258 23828 16270
rect 23884 16212 23940 16222
rect 23884 16118 23940 16156
rect 23212 15934 23214 15986
rect 23266 15934 23268 15986
rect 23212 15922 23268 15934
rect 22540 15374 22542 15426
rect 22594 15374 22596 15426
rect 22540 15362 22596 15374
rect 21868 15262 21870 15314
rect 21922 15262 21924 15314
rect 21868 15250 21924 15262
rect 23996 15204 24052 16828
rect 24556 16818 24612 16828
rect 24668 15204 24724 15214
rect 23996 15202 24724 15204
rect 23996 15150 24670 15202
rect 24722 15150 24724 15202
rect 23996 15148 24724 15150
rect 19628 14578 19684 14588
rect 20636 14642 20804 14644
rect 20636 14590 20750 14642
rect 20802 14590 20804 14642
rect 20636 14588 20804 14590
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20300 13634 20356 13646
rect 20300 13582 20302 13634
rect 20354 13582 20356 13634
rect 20300 13524 20356 13582
rect 20300 13458 20356 13468
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19516 8372 19684 8428
rect 19628 4340 19684 8372
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19740 4340 19796 4350
rect 19628 4338 19796 4340
rect 19628 4286 19742 4338
rect 19794 4286 19796 4338
rect 19628 4284 19796 4286
rect 19740 4274 19796 4284
rect 19852 4116 19908 4126
rect 19740 3556 19796 3566
rect 19404 3554 19796 3556
rect 19404 3502 19742 3554
rect 19794 3502 19796 3554
rect 19404 3500 19796 3502
rect 19740 3490 19796 3500
rect 19852 3332 19908 4060
rect 20636 3556 20692 14588
rect 20748 14578 20804 14588
rect 20748 13748 20804 13758
rect 20748 13654 20804 13692
rect 24668 13524 24724 15148
rect 24444 13468 24724 13524
rect 24444 8428 24500 13468
rect 24780 8428 24836 17164
rect 25676 16098 25732 17948
rect 25788 17108 25844 17118
rect 25788 16882 25844 17052
rect 25788 16830 25790 16882
rect 25842 16830 25844 16882
rect 25788 16818 25844 16830
rect 25676 16046 25678 16098
rect 25730 16046 25732 16098
rect 25340 15316 25396 15326
rect 25676 15316 25732 16046
rect 26012 16770 26068 16782
rect 26012 16718 26014 16770
rect 26066 16718 26068 16770
rect 26012 15426 26068 16718
rect 26348 16772 26404 18510
rect 26460 18676 26516 18686
rect 26460 18450 26516 18620
rect 27020 18564 27076 22428
rect 27132 21588 27188 23102
rect 27356 22260 27412 23212
rect 28364 23268 28420 23774
rect 28364 23202 28420 23212
rect 30044 23380 30100 23390
rect 27916 23044 27972 23054
rect 30044 23044 30100 23324
rect 37660 23380 37716 23886
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 37660 23314 37716 23324
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 27916 23042 28532 23044
rect 27916 22990 27918 23042
rect 27970 22990 28532 23042
rect 27916 22988 28532 22990
rect 27916 22978 27972 22988
rect 28476 22594 28532 22988
rect 29484 23042 30100 23044
rect 29484 22990 30046 23042
rect 30098 22990 30100 23042
rect 29484 22988 30100 22990
rect 28476 22542 28478 22594
rect 28530 22542 28532 22594
rect 28476 22530 28532 22542
rect 28812 22540 29316 22596
rect 28588 22484 28644 22494
rect 28812 22484 28868 22540
rect 28588 22482 28868 22484
rect 28588 22430 28590 22482
rect 28642 22430 28868 22482
rect 28588 22428 28868 22430
rect 29260 22482 29316 22540
rect 29260 22430 29262 22482
rect 29314 22430 29316 22482
rect 28588 22418 28644 22428
rect 29260 22418 29316 22430
rect 27356 22166 27412 22204
rect 27468 22372 27524 22382
rect 27468 22258 27524 22316
rect 27692 22372 27748 22382
rect 28140 22372 28196 22382
rect 27692 22370 28196 22372
rect 27692 22318 27694 22370
rect 27746 22318 28142 22370
rect 28194 22318 28196 22370
rect 27692 22316 28196 22318
rect 27692 22306 27748 22316
rect 28140 22306 28196 22316
rect 29036 22370 29092 22382
rect 29036 22318 29038 22370
rect 29090 22318 29092 22370
rect 27468 22206 27470 22258
rect 27522 22206 27524 22258
rect 27468 22194 27524 22206
rect 29036 22260 29092 22318
rect 29484 22370 29540 22988
rect 30044 22978 30100 22988
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 29484 22318 29486 22370
rect 29538 22318 29540 22370
rect 29484 22306 29540 22318
rect 29596 22484 29652 22494
rect 29596 22370 29652 22428
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 29596 22318 29598 22370
rect 29650 22318 29652 22370
rect 29596 22306 29652 22318
rect 30044 22372 30100 22382
rect 29036 22194 29092 22204
rect 27804 22146 27860 22158
rect 27804 22094 27806 22146
rect 27858 22094 27860 22146
rect 27804 21700 27860 22094
rect 28028 22146 28084 22158
rect 28028 22094 28030 22146
rect 28082 22094 28084 22146
rect 27916 21700 27972 21710
rect 27804 21698 27972 21700
rect 27804 21646 27918 21698
rect 27970 21646 27972 21698
rect 27804 21644 27972 21646
rect 27916 21634 27972 21644
rect 27132 21494 27188 21532
rect 28028 21140 28084 22094
rect 30044 21474 30100 22316
rect 37660 22372 37716 22382
rect 37660 22278 37716 22316
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 30044 21422 30046 21474
rect 30098 21422 30100 21474
rect 30044 21410 30100 21422
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 27356 21084 28084 21140
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 27356 19234 27412 21084
rect 27468 20916 27524 20926
rect 27468 20020 27524 20860
rect 28588 20132 28644 20142
rect 27468 20018 28084 20020
rect 27468 19966 27470 20018
rect 27522 19966 28084 20018
rect 27468 19964 28084 19966
rect 27468 19954 27524 19964
rect 27468 19348 27524 19358
rect 27468 19346 27972 19348
rect 27468 19294 27470 19346
rect 27522 19294 27972 19346
rect 27468 19292 27972 19294
rect 27468 19282 27524 19292
rect 27356 19182 27358 19234
rect 27410 19182 27412 19234
rect 27132 19012 27188 19022
rect 27132 18918 27188 18956
rect 27356 18674 27412 19182
rect 27916 19234 27972 19292
rect 27916 19182 27918 19234
rect 27970 19182 27972 19234
rect 27916 19170 27972 19182
rect 27356 18622 27358 18674
rect 27410 18622 27412 18674
rect 27356 18610 27412 18622
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 26460 18386 26516 18398
rect 26908 18562 27076 18564
rect 26908 18510 27022 18562
rect 27074 18510 27076 18562
rect 26908 18508 27076 18510
rect 26908 17220 26964 18508
rect 27020 18498 27076 18508
rect 27132 18564 27188 18574
rect 27132 18562 27300 18564
rect 27132 18510 27134 18562
rect 27186 18510 27300 18562
rect 27132 18508 27300 18510
rect 27132 18498 27188 18508
rect 26852 17164 26964 17220
rect 26460 16996 26516 17006
rect 26460 16902 26516 16940
rect 26684 16884 26740 16894
rect 26852 16884 26908 17164
rect 27244 16996 27300 18508
rect 27804 18452 27860 18462
rect 28028 18452 28084 19964
rect 28252 19908 28308 19918
rect 28252 19814 28308 19852
rect 28588 19236 28644 20076
rect 30716 20020 30772 20030
rect 29484 19908 29540 19918
rect 30380 19908 30436 19918
rect 28588 19142 28644 19180
rect 29260 19236 29316 19246
rect 29260 19142 29316 19180
rect 28364 19122 28420 19134
rect 28364 19070 28366 19122
rect 28418 19070 28420 19122
rect 28252 19010 28308 19022
rect 28252 18958 28254 19010
rect 28306 18958 28308 19010
rect 28252 18676 28308 18958
rect 28364 19012 28420 19070
rect 28364 18946 28420 18956
rect 29372 19122 29428 19134
rect 29372 19070 29374 19122
rect 29426 19070 29428 19122
rect 29372 18676 29428 19070
rect 29484 19010 29540 19852
rect 30156 19906 30436 19908
rect 30156 19854 30382 19906
rect 30434 19854 30436 19906
rect 30156 19852 30436 19854
rect 30156 19236 30212 19852
rect 30380 19842 30436 19852
rect 29708 19124 29764 19134
rect 29932 19124 29988 19134
rect 29708 19122 29988 19124
rect 29708 19070 29710 19122
rect 29762 19070 29934 19122
rect 29986 19070 29988 19122
rect 29708 19068 29988 19070
rect 29708 19058 29764 19068
rect 29932 19058 29988 19068
rect 30156 19122 30212 19180
rect 30156 19070 30158 19122
rect 30210 19070 30212 19122
rect 30156 19058 30212 19070
rect 30268 19124 30324 19134
rect 30604 19124 30660 19134
rect 30268 19122 30660 19124
rect 30268 19070 30270 19122
rect 30322 19070 30606 19122
rect 30658 19070 30660 19122
rect 30268 19068 30660 19070
rect 29484 18958 29486 19010
rect 29538 18958 29540 19010
rect 29484 18946 29540 18958
rect 28252 18620 28532 18676
rect 28476 18562 28532 18620
rect 29372 18610 29428 18620
rect 28476 18510 28478 18562
rect 28530 18510 28532 18562
rect 28476 18498 28532 18510
rect 27804 18450 28084 18452
rect 27804 18398 27806 18450
rect 27858 18398 28084 18450
rect 27804 18396 28084 18398
rect 27804 18004 27860 18396
rect 27804 17938 27860 17948
rect 27244 16930 27300 16940
rect 27356 17164 28420 17220
rect 27356 16994 27412 17164
rect 28364 17106 28420 17164
rect 28364 17054 28366 17106
rect 28418 17054 28420 17106
rect 28364 17042 28420 17054
rect 27356 16942 27358 16994
rect 27410 16942 27412 16994
rect 27356 16930 27412 16942
rect 30268 16996 30324 19068
rect 30604 19058 30660 19068
rect 30716 19122 30772 19964
rect 37660 20020 37716 20030
rect 37660 19926 37716 19964
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37884 19348 37940 21534
rect 40012 21362 40068 21374
rect 40012 21310 40014 21362
rect 40066 21310 40068 21362
rect 40012 20916 40068 21310
rect 40012 20850 40068 20860
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37884 19282 37940 19292
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 30716 19070 30718 19122
rect 30770 19070 30772 19122
rect 30604 18340 30660 18350
rect 30716 18340 30772 19070
rect 30940 19012 30996 19022
rect 30940 18918 30996 18956
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 30604 18338 30772 18340
rect 30604 18286 30606 18338
rect 30658 18286 30772 18338
rect 30604 18284 30772 18286
rect 30604 18274 30660 18284
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 30268 16930 30324 16940
rect 26684 16882 26908 16884
rect 26684 16830 26686 16882
rect 26738 16830 26908 16882
rect 26684 16828 26908 16830
rect 27132 16884 27188 16894
rect 26684 16818 26740 16828
rect 27132 16790 27188 16828
rect 28028 16882 28084 16894
rect 28028 16830 28030 16882
rect 28082 16830 28084 16882
rect 26124 16660 26180 16670
rect 26124 16566 26180 16604
rect 26348 16212 26404 16716
rect 26572 16770 26628 16782
rect 26572 16718 26574 16770
rect 26626 16718 26628 16770
rect 26348 16146 26404 16156
rect 26460 16212 26516 16222
rect 26572 16212 26628 16718
rect 27468 16772 27524 16782
rect 27692 16772 27748 16782
rect 27524 16770 27748 16772
rect 27524 16718 27694 16770
rect 27746 16718 27748 16770
rect 27524 16716 27748 16718
rect 27468 16706 27524 16716
rect 27692 16706 27748 16716
rect 27804 16772 27860 16782
rect 27804 16678 27860 16716
rect 26908 16658 26964 16670
rect 26908 16606 26910 16658
rect 26962 16606 26964 16658
rect 26908 16548 26964 16606
rect 26908 16482 26964 16492
rect 26460 16210 26628 16212
rect 26460 16158 26462 16210
rect 26514 16158 26628 16210
rect 26460 16156 26628 16158
rect 26460 16146 26516 16156
rect 28028 16100 28084 16830
rect 28476 16884 28532 16894
rect 37660 16884 37716 16894
rect 28532 16828 28644 16884
rect 28476 16790 28532 16828
rect 28588 16210 28644 16828
rect 37660 16790 37716 16828
rect 39900 16770 39956 16782
rect 39900 16718 39902 16770
rect 39954 16718 39956 16770
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 28588 16158 28590 16210
rect 28642 16158 28644 16210
rect 28588 16146 28644 16158
rect 39900 16212 39956 16718
rect 39900 16146 39956 16156
rect 40012 16210 40068 16222
rect 40012 16158 40014 16210
rect 40066 16158 40068 16210
rect 37660 16100 37716 16110
rect 28084 16044 28196 16100
rect 28028 16034 28084 16044
rect 26012 15374 26014 15426
rect 26066 15374 26068 15426
rect 26012 15362 26068 15374
rect 25340 15314 25732 15316
rect 25340 15262 25342 15314
rect 25394 15262 25732 15314
rect 25340 15260 25732 15262
rect 25340 15250 25396 15260
rect 28140 15202 28196 16044
rect 37660 16006 37716 16044
rect 40012 15540 40068 16158
rect 40012 15474 40068 15484
rect 28140 15150 28142 15202
rect 28194 15150 28196 15202
rect 28140 15138 28196 15150
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 23772 8372 24500 8428
rect 24556 8372 24836 8428
rect 23548 5236 23604 5246
rect 20748 4116 20804 4126
rect 20748 4022 20804 4060
rect 22876 3668 22932 3678
rect 20748 3556 20804 3566
rect 20636 3554 20804 3556
rect 20636 3502 20750 3554
rect 20802 3502 20804 3554
rect 20636 3500 20804 3502
rect 20748 3490 20804 3500
rect 19516 3276 19908 3332
rect 20188 3444 20244 3454
rect 19516 800 19572 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 3388
rect 21756 3444 21812 3454
rect 21756 3330 21812 3388
rect 21756 3278 21758 3330
rect 21810 3278 21812 3330
rect 21756 3266 21812 3278
rect 22876 800 22932 3612
rect 23548 800 23604 5180
rect 23772 5122 23828 8372
rect 23772 5070 23774 5122
rect 23826 5070 23828 5122
rect 23772 5058 23828 5070
rect 24556 3554 24612 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 24780 5236 24836 5246
rect 24780 5142 24836 5180
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 35980 3332 36036 3342
rect 35644 3330 36036 3332
rect 35644 3278 35982 3330
rect 36034 3278 36036 3330
rect 35644 3276 36036 3278
rect 35644 800 35700 3276
rect 35980 3266 36036 3276
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 35616 0 35728 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 15484 36652 15540 36708
rect 16716 36706 16772 36708
rect 16716 36654 16718 36706
rect 16718 36654 16770 36706
rect 16770 36654 16772 36706
rect 16716 36652 16772 36654
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 27580 4228 27636
rect 1932 26236 1988 26292
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 11788 27020 11844 27076
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 13356 26908 13412 26964
rect 14252 26962 14308 26964
rect 14252 26910 14254 26962
rect 14254 26910 14306 26962
rect 14306 26910 14308 26962
rect 14252 26908 14308 26910
rect 11788 25452 11844 25508
rect 14364 26236 14420 26292
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 25564 38556 25620 38612
rect 26796 38556 26852 38612
rect 24892 38220 24948 38276
rect 26124 38274 26180 38276
rect 26124 38222 26126 38274
rect 26126 38222 26178 38274
rect 26178 38222 26180 38274
rect 26124 38220 26180 38222
rect 21532 37436 21588 37492
rect 22764 37490 22820 37492
rect 22764 37438 22766 37490
rect 22766 37438 22818 37490
rect 22818 37438 22820 37490
rect 22764 37436 22820 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19516 28476 19572 28532
rect 17612 27804 17668 27860
rect 18172 27804 18228 27860
rect 14924 25900 14980 25956
rect 14700 25506 14756 25508
rect 14700 25454 14702 25506
rect 14702 25454 14754 25506
rect 14754 25454 14756 25506
rect 14700 25452 14756 25454
rect 17388 26908 17444 26964
rect 15820 26124 15876 26180
rect 15372 25228 15428 25284
rect 12684 24668 12740 24724
rect 14588 24722 14644 24724
rect 14588 24670 14590 24722
rect 14590 24670 14642 24722
rect 14642 24670 14644 24722
rect 14588 24668 14644 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 12012 23324 12068 23380
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 21420 4228 21476
rect 14140 22540 14196 22596
rect 14140 22316 14196 22372
rect 12124 22092 12180 22148
rect 13916 22146 13972 22148
rect 13916 22094 13918 22146
rect 13918 22094 13970 22146
rect 13970 22094 13972 22146
rect 13916 22092 13972 22094
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 14924 22540 14980 22596
rect 14924 22092 14980 22148
rect 15148 24722 15204 24724
rect 15148 24670 15150 24722
rect 15150 24670 15202 24722
rect 15202 24670 15204 24722
rect 15148 24668 15204 24670
rect 15932 25900 15988 25956
rect 16156 26290 16212 26292
rect 16156 26238 16158 26290
rect 16158 26238 16210 26290
rect 16210 26238 16212 26290
rect 16156 26236 16212 26238
rect 17388 26124 17444 26180
rect 16380 25452 16436 25508
rect 16268 25394 16324 25396
rect 16268 25342 16270 25394
rect 16270 25342 16322 25394
rect 16322 25342 16324 25394
rect 16268 25340 16324 25342
rect 17500 25506 17556 25508
rect 17500 25454 17502 25506
rect 17502 25454 17554 25506
rect 17554 25454 17556 25506
rect 17500 25452 17556 25454
rect 16380 25228 16436 25284
rect 15708 24668 15764 24724
rect 17276 25228 17332 25284
rect 17948 25506 18004 25508
rect 17948 25454 17950 25506
rect 17950 25454 18002 25506
rect 18002 25454 18004 25506
rect 17948 25452 18004 25454
rect 19068 27468 19124 27524
rect 18844 26908 18900 26964
rect 20972 28476 21028 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 22540 28082 22596 28084
rect 22540 28030 22542 28082
rect 22542 28030 22594 28082
rect 22594 28030 22596 28082
rect 22540 28028 22596 28030
rect 19516 27020 19572 27076
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 23548 28028 23604 28084
rect 19964 26908 20020 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20188 26460 20244 26516
rect 20300 26796 20356 26852
rect 19628 26348 19684 26404
rect 20860 26796 20916 26852
rect 22204 26796 22260 26852
rect 22428 26908 22484 26964
rect 21420 26514 21476 26516
rect 21420 26462 21422 26514
rect 21422 26462 21474 26514
rect 21474 26462 21476 26514
rect 21420 26460 21476 26462
rect 16492 24668 16548 24724
rect 18508 24498 18564 24500
rect 18508 24446 18510 24498
rect 18510 24446 18562 24498
rect 18562 24446 18564 24498
rect 18508 24444 18564 24446
rect 18732 24722 18788 24724
rect 18732 24670 18734 24722
rect 18734 24670 18786 24722
rect 18786 24670 18788 24722
rect 18732 24668 18788 24670
rect 15260 23212 15316 23268
rect 17388 23266 17444 23268
rect 17388 23214 17390 23266
rect 17390 23214 17442 23266
rect 17442 23214 17444 23266
rect 17388 23212 17444 23214
rect 17724 23154 17780 23156
rect 17724 23102 17726 23154
rect 17726 23102 17778 23154
rect 17778 23102 17780 23154
rect 17724 23100 17780 23102
rect 16380 22482 16436 22484
rect 16380 22430 16382 22482
rect 16382 22430 16434 22482
rect 16434 22430 16436 22482
rect 16380 22428 16436 22430
rect 15372 22316 15428 22372
rect 16156 22370 16212 22372
rect 16156 22318 16158 22370
rect 16158 22318 16210 22370
rect 16210 22318 16212 22370
rect 16156 22316 16212 22318
rect 17388 22370 17444 22372
rect 17388 22318 17390 22370
rect 17390 22318 17442 22370
rect 17442 22318 17444 22370
rect 17388 22316 17444 22318
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 14140 19964 14196 20020
rect 12012 19906 12068 19908
rect 12012 19854 12014 19906
rect 12014 19854 12066 19906
rect 12066 19854 12068 19906
rect 12012 19852 12068 19854
rect 14476 19906 14532 19908
rect 14476 19854 14478 19906
rect 14478 19854 14530 19906
rect 14530 19854 14532 19906
rect 14476 19852 14532 19854
rect 14588 19404 14644 19460
rect 11340 18956 11396 19012
rect 13804 19010 13860 19012
rect 13804 18958 13806 19010
rect 13806 18958 13858 19010
rect 13858 18958 13860 19010
rect 13804 18956 13860 18958
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 10668 18396 10724 18452
rect 14028 18844 14084 18900
rect 12348 18284 12404 18340
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 14252 18396 14308 18452
rect 15148 20914 15204 20916
rect 15148 20862 15150 20914
rect 15150 20862 15202 20914
rect 15202 20862 15204 20914
rect 15148 20860 15204 20862
rect 15484 20636 15540 20692
rect 18172 22428 18228 22484
rect 18956 25452 19012 25508
rect 20524 26348 20580 26404
rect 20076 25394 20132 25396
rect 20076 25342 20078 25394
rect 20078 25342 20130 25394
rect 20130 25342 20132 25394
rect 20076 25340 20132 25342
rect 19180 25228 19236 25284
rect 18956 24892 19012 24948
rect 19180 24668 19236 24724
rect 18956 24444 19012 24500
rect 18620 23212 18676 23268
rect 18956 23212 19012 23268
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19628 24332 19684 24388
rect 20188 24332 20244 24388
rect 20300 25340 20356 25396
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20748 26402 20804 26404
rect 20748 26350 20750 26402
rect 20750 26350 20802 26402
rect 20802 26350 20804 26402
rect 20748 26348 20804 26350
rect 22540 26236 22596 26292
rect 22316 25564 22372 25620
rect 22428 25394 22484 25396
rect 22428 25342 22430 25394
rect 22430 25342 22482 25394
rect 22482 25342 22484 25394
rect 22428 25340 22484 25342
rect 22316 25228 22372 25284
rect 22540 25228 22596 25284
rect 22652 25900 22708 25956
rect 20524 24892 20580 24948
rect 20748 24722 20804 24724
rect 20748 24670 20750 24722
rect 20750 24670 20802 24722
rect 20802 24670 20804 24722
rect 20748 24668 20804 24670
rect 20300 23324 20356 23380
rect 20860 23378 20916 23380
rect 20860 23326 20862 23378
rect 20862 23326 20914 23378
rect 20914 23326 20916 23378
rect 20860 23324 20916 23326
rect 19068 23154 19124 23156
rect 19068 23102 19070 23154
rect 19070 23102 19122 23154
rect 19122 23102 19124 23154
rect 19068 23100 19124 23102
rect 18732 22988 18788 23044
rect 19964 23100 20020 23156
rect 20636 23154 20692 23156
rect 20636 23102 20638 23154
rect 20638 23102 20690 23154
rect 20690 23102 20692 23154
rect 20636 23100 20692 23102
rect 18620 22540 18676 22596
rect 19628 22988 19684 23044
rect 18508 22316 18564 22372
rect 17836 21868 17892 21924
rect 18284 21868 18340 21924
rect 17500 21698 17556 21700
rect 17500 21646 17502 21698
rect 17502 21646 17554 21698
rect 17554 21646 17556 21698
rect 17500 21644 17556 21646
rect 17948 21644 18004 21700
rect 16828 21474 16884 21476
rect 16828 21422 16830 21474
rect 16830 21422 16882 21474
rect 16882 21422 16884 21474
rect 16828 21420 16884 21422
rect 14700 18956 14756 19012
rect 15260 20018 15316 20020
rect 15260 19966 15262 20018
rect 15262 19966 15314 20018
rect 15314 19966 15316 20018
rect 15260 19964 15316 19966
rect 15596 19628 15652 19684
rect 15932 19404 15988 19460
rect 16044 19628 16100 19684
rect 14588 18844 14644 18900
rect 14700 18732 14756 18788
rect 14476 18508 14532 18564
rect 14140 18338 14196 18340
rect 14140 18286 14142 18338
rect 14142 18286 14194 18338
rect 14194 18286 14196 18338
rect 14140 18284 14196 18286
rect 14252 16940 14308 16996
rect 4284 16882 4340 16884
rect 4284 16830 4286 16882
rect 4286 16830 4338 16882
rect 4338 16830 4340 16882
rect 4284 16828 4340 16830
rect 12460 16828 12516 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 16156 1988 16212
rect 16492 19068 16548 19124
rect 17052 19122 17108 19124
rect 17052 19070 17054 19122
rect 17054 19070 17106 19122
rect 17106 19070 17108 19122
rect 17052 19068 17108 19070
rect 15372 19010 15428 19012
rect 15372 18958 15374 19010
rect 15374 18958 15426 19010
rect 15426 18958 15428 19010
rect 15372 18956 15428 18958
rect 15260 18620 15316 18676
rect 15036 16994 15092 16996
rect 15036 16942 15038 16994
rect 15038 16942 15090 16994
rect 15090 16942 15092 16994
rect 15036 16940 15092 16942
rect 16716 18620 16772 18676
rect 15708 18508 15764 18564
rect 14924 16604 14980 16660
rect 15372 16828 15428 16884
rect 12460 15932 12516 15988
rect 16828 18338 16884 18340
rect 16828 18286 16830 18338
rect 16830 18286 16882 18338
rect 16882 18286 16884 18338
rect 16828 18284 16884 18286
rect 16380 17612 16436 17668
rect 17388 19068 17444 19124
rect 17836 20300 17892 20356
rect 17948 20860 18004 20916
rect 17612 19068 17668 19124
rect 17948 19068 18004 19124
rect 17500 18956 17556 19012
rect 17836 18956 17892 19012
rect 15708 16828 15764 16884
rect 16828 17388 16884 17444
rect 17724 18732 17780 18788
rect 17948 18732 18004 18788
rect 17948 18396 18004 18452
rect 17724 17666 17780 17668
rect 17724 17614 17726 17666
rect 17726 17614 17778 17666
rect 17778 17614 17780 17666
rect 17724 17612 17780 17614
rect 17164 16940 17220 16996
rect 17388 16882 17444 16884
rect 17388 16830 17390 16882
rect 17390 16830 17442 16882
rect 17442 16830 17444 16882
rect 17388 16828 17444 16830
rect 15484 16716 15540 16772
rect 16268 16716 16324 16772
rect 15820 16492 15876 16548
rect 15596 15986 15652 15988
rect 15596 15934 15598 15986
rect 15598 15934 15650 15986
rect 15650 15934 15652 15986
rect 15596 15932 15652 15934
rect 14028 15148 14084 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 16604 16770 16660 16772
rect 16604 16718 16606 16770
rect 16606 16718 16658 16770
rect 16658 16718 16660 16770
rect 16604 16716 16660 16718
rect 17276 16716 17332 16772
rect 16492 16658 16548 16660
rect 16492 16606 16494 16658
rect 16494 16606 16546 16658
rect 16546 16606 16548 16658
rect 16492 16604 16548 16606
rect 18956 22482 19012 22484
rect 18956 22430 18958 22482
rect 18958 22430 19010 22482
rect 19010 22430 19012 22482
rect 18956 22428 19012 22430
rect 19516 22428 19572 22484
rect 19068 22316 19124 22372
rect 18732 20188 18788 20244
rect 19292 22316 19348 22372
rect 19180 21868 19236 21924
rect 19068 20188 19124 20244
rect 18620 19628 18676 19684
rect 18732 19794 18788 19796
rect 18732 19742 18734 19794
rect 18734 19742 18786 19794
rect 18786 19742 18788 19794
rect 18732 19740 18788 19742
rect 18508 18620 18564 18676
rect 18620 18450 18676 18452
rect 18620 18398 18622 18450
rect 18622 18398 18674 18450
rect 18674 18398 18676 18450
rect 18620 18396 18676 18398
rect 18172 18284 18228 18340
rect 18508 18284 18564 18340
rect 18060 17836 18116 17892
rect 18396 17442 18452 17444
rect 18396 17390 18398 17442
rect 18398 17390 18450 17442
rect 18450 17390 18452 17442
rect 18396 17388 18452 17390
rect 17612 16492 17668 16548
rect 15708 15202 15764 15204
rect 15708 15150 15710 15202
rect 15710 15150 15762 15202
rect 15762 15150 15764 15202
rect 15708 15148 15764 15150
rect 17612 15148 17668 15204
rect 18060 16828 18116 16884
rect 18284 16492 18340 16548
rect 15596 14306 15652 14308
rect 15596 14254 15598 14306
rect 15598 14254 15650 14306
rect 15650 14254 15652 14306
rect 15596 14252 15652 14254
rect 17500 14306 17556 14308
rect 17500 14254 17502 14306
rect 17502 14254 17554 14306
rect 17554 14254 17556 14306
rect 17500 14252 17556 14254
rect 19404 21420 19460 21476
rect 19404 20300 19460 20356
rect 19180 19964 19236 20020
rect 19404 18450 19460 18452
rect 19404 18398 19406 18450
rect 19406 18398 19458 18450
rect 19458 18398 19460 18450
rect 19404 18396 19460 18398
rect 19292 18284 19348 18340
rect 18956 17612 19012 17668
rect 19068 17836 19124 17892
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 22316 24722 22372 24724
rect 22316 24670 22318 24722
rect 22318 24670 22370 24722
rect 22370 24670 22372 24722
rect 22316 24668 22372 24670
rect 23660 26908 23716 26964
rect 23884 26514 23940 26516
rect 23884 26462 23886 26514
rect 23886 26462 23938 26514
rect 23938 26462 23940 26514
rect 23884 26460 23940 26462
rect 22988 26178 23044 26180
rect 22988 26126 22990 26178
rect 22990 26126 23042 26178
rect 23042 26126 23044 26178
rect 22988 26124 23044 26126
rect 23100 26066 23156 26068
rect 23100 26014 23102 26066
rect 23102 26014 23154 26066
rect 23154 26014 23156 26066
rect 23100 26012 23156 26014
rect 23660 26290 23716 26292
rect 23660 26238 23662 26290
rect 23662 26238 23714 26290
rect 23714 26238 23716 26290
rect 23660 26236 23716 26238
rect 23996 26290 24052 26292
rect 23996 26238 23998 26290
rect 23998 26238 24050 26290
rect 24050 26238 24052 26290
rect 23996 26236 24052 26238
rect 23772 26178 23828 26180
rect 23772 26126 23774 26178
rect 23774 26126 23826 26178
rect 23826 26126 23828 26178
rect 23772 26124 23828 26126
rect 23324 25564 23380 25620
rect 21308 22482 21364 22484
rect 21308 22430 21310 22482
rect 21310 22430 21362 22482
rect 21362 22430 21364 22482
rect 21308 22428 21364 22430
rect 22652 23436 22708 23492
rect 20636 22204 20692 22260
rect 21644 22258 21700 22260
rect 21644 22206 21646 22258
rect 21646 22206 21698 22258
rect 21698 22206 21700 22258
rect 21644 22204 21700 22206
rect 20076 21644 20132 21700
rect 20076 21420 20132 21476
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 21420 20188 21476 20244
rect 21532 20636 21588 20692
rect 19740 19740 19796 19796
rect 20412 19964 20468 20020
rect 20300 19628 20356 19684
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 21308 20018 21364 20020
rect 21308 19966 21310 20018
rect 21310 19966 21362 20018
rect 21362 19966 21364 20018
rect 21308 19964 21364 19966
rect 22652 22258 22708 22260
rect 22652 22206 22654 22258
rect 22654 22206 22706 22258
rect 22706 22206 22708 22258
rect 22652 22204 22708 22206
rect 22652 21026 22708 21028
rect 22652 20974 22654 21026
rect 22654 20974 22706 21026
rect 22706 20974 22708 21026
rect 22652 20972 22708 20974
rect 22764 20860 22820 20916
rect 22652 20802 22708 20804
rect 22652 20750 22654 20802
rect 22654 20750 22706 20802
rect 22706 20750 22708 20802
rect 22652 20748 22708 20750
rect 22316 20690 22372 20692
rect 22316 20638 22318 20690
rect 22318 20638 22370 20690
rect 22370 20638 22372 20690
rect 22316 20636 22372 20638
rect 21644 19628 21700 19684
rect 21756 19458 21812 19460
rect 21756 19406 21758 19458
rect 21758 19406 21810 19458
rect 21810 19406 21812 19458
rect 21756 19404 21812 19406
rect 22316 18956 22372 19012
rect 20860 18396 20916 18452
rect 19628 17836 19684 17892
rect 19628 17554 19684 17556
rect 19628 17502 19630 17554
rect 19630 17502 19682 17554
rect 19682 17502 19684 17554
rect 19628 17500 19684 17502
rect 18732 17164 18788 17220
rect 18732 16828 18788 16884
rect 19628 17276 19684 17332
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19740 16828 19796 16884
rect 20076 16604 20132 16660
rect 18732 15484 18788 15540
rect 17500 13746 17556 13748
rect 17500 13694 17502 13746
rect 17502 13694 17554 13746
rect 17554 13694 17556 13746
rect 17500 13692 17556 13694
rect 18732 14588 18788 14644
rect 18508 13468 18564 13524
rect 19404 13468 19460 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 22204 17836 22260 17892
rect 21868 17612 21924 17668
rect 20860 17500 20916 17556
rect 21420 17106 21476 17108
rect 21420 17054 21422 17106
rect 21422 17054 21474 17106
rect 21474 17054 21476 17106
rect 21420 17052 21476 17054
rect 21084 16658 21140 16660
rect 21084 16606 21086 16658
rect 21086 16606 21138 16658
rect 21138 16606 21140 16658
rect 21084 16604 21140 16606
rect 20412 16156 20468 16212
rect 20524 15202 20580 15204
rect 20524 15150 20526 15202
rect 20526 15150 20578 15202
rect 20578 15150 20580 15202
rect 20524 15148 20580 15150
rect 22876 17612 22932 17668
rect 22988 20076 23044 20132
rect 23660 26012 23716 26068
rect 24556 27132 24612 27188
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 25900 27186 25956 27188
rect 25900 27134 25902 27186
rect 25902 27134 25954 27186
rect 25954 27134 25956 27186
rect 25900 27132 25956 27134
rect 25788 26460 25844 26516
rect 24444 26290 24500 26292
rect 24444 26238 24446 26290
rect 24446 26238 24498 26290
rect 24498 26238 24500 26290
rect 24444 26236 24500 26238
rect 23996 25900 24052 25956
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 23436 25228 23492 25284
rect 25900 24332 25956 24388
rect 25900 23660 25956 23716
rect 24556 23436 24612 23492
rect 24444 22876 24500 22932
rect 23212 20972 23268 21028
rect 23324 21474 23380 21476
rect 23324 21422 23326 21474
rect 23326 21422 23378 21474
rect 23378 21422 23380 21474
rect 23324 21420 23380 21422
rect 23100 18956 23156 19012
rect 23884 21196 23940 21252
rect 24668 22876 24724 22932
rect 24780 22258 24836 22260
rect 24780 22206 24782 22258
rect 24782 22206 24834 22258
rect 24834 22206 24836 22258
rect 24780 22204 24836 22206
rect 24220 20748 24276 20804
rect 25228 21196 25284 21252
rect 23772 20130 23828 20132
rect 23772 20078 23774 20130
rect 23774 20078 23826 20130
rect 23826 20078 23828 20130
rect 23772 20076 23828 20078
rect 22652 17164 22708 17220
rect 22764 16994 22820 16996
rect 22764 16942 22766 16994
rect 22766 16942 22818 16994
rect 22818 16942 22820 16994
rect 22764 16940 22820 16942
rect 22428 16882 22484 16884
rect 22428 16830 22430 16882
rect 22430 16830 22482 16882
rect 22482 16830 22484 16882
rect 22428 16828 22484 16830
rect 23324 18450 23380 18452
rect 23324 18398 23326 18450
rect 23326 18398 23378 18450
rect 23378 18398 23380 18450
rect 23324 18396 23380 18398
rect 23212 16882 23268 16884
rect 23212 16830 23214 16882
rect 23214 16830 23266 16882
rect 23266 16830 23268 16882
rect 23212 16828 23268 16830
rect 25340 20914 25396 20916
rect 25340 20862 25342 20914
rect 25342 20862 25394 20914
rect 25394 20862 25396 20914
rect 25340 20860 25396 20862
rect 25788 19346 25844 19348
rect 25788 19294 25790 19346
rect 25790 19294 25842 19346
rect 25842 19294 25844 19346
rect 25788 19292 25844 19294
rect 28252 24668 28308 24724
rect 29484 24668 29540 24724
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 27468 23714 27524 23716
rect 27468 23662 27470 23714
rect 27470 23662 27522 23714
rect 27522 23662 27524 23714
rect 27468 23660 27524 23662
rect 27356 23212 27412 23268
rect 26572 21532 26628 21588
rect 26572 20860 26628 20916
rect 27020 22428 27076 22484
rect 26124 18956 26180 19012
rect 26908 19010 26964 19012
rect 26908 18958 26910 19010
rect 26910 18958 26962 19010
rect 26962 18958 26964 19010
rect 26908 18956 26964 18958
rect 26348 18732 26404 18788
rect 25676 17948 25732 18004
rect 24556 17164 24612 17220
rect 23884 16210 23940 16212
rect 23884 16158 23886 16210
rect 23886 16158 23938 16210
rect 23938 16158 23940 16210
rect 23884 16156 23940 16158
rect 24556 16828 24612 16884
rect 19628 14588 19684 14644
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20300 13468 20356 13524
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19852 4060 19908 4116
rect 20748 13746 20804 13748
rect 20748 13694 20750 13746
rect 20750 13694 20802 13746
rect 20802 13694 20804 13746
rect 20748 13692 20804 13694
rect 25788 17052 25844 17108
rect 26460 18620 26516 18676
rect 28364 23212 28420 23268
rect 30044 23324 30100 23380
rect 40012 23548 40068 23604
rect 37660 23324 37716 23380
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 27356 22258 27412 22260
rect 27356 22206 27358 22258
rect 27358 22206 27410 22258
rect 27410 22206 27412 22258
rect 27356 22204 27412 22206
rect 27468 22316 27524 22372
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 29596 22428 29652 22484
rect 30044 22316 30100 22372
rect 29036 22204 29092 22260
rect 27132 21586 27188 21588
rect 27132 21534 27134 21586
rect 27134 21534 27186 21586
rect 27186 21534 27188 21586
rect 27132 21532 27188 21534
rect 37660 22370 37716 22372
rect 37660 22318 37662 22370
rect 37662 22318 37714 22370
rect 37714 22318 37716 22370
rect 37660 22316 37716 22318
rect 40012 22204 40068 22260
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 27468 20860 27524 20916
rect 28588 20076 28644 20132
rect 27132 19010 27188 19012
rect 27132 18958 27134 19010
rect 27134 18958 27186 19010
rect 27186 18958 27188 19010
rect 27132 18956 27188 18958
rect 26460 16994 26516 16996
rect 26460 16942 26462 16994
rect 26462 16942 26514 16994
rect 26514 16942 26516 16994
rect 26460 16940 26516 16942
rect 28252 19906 28308 19908
rect 28252 19854 28254 19906
rect 28254 19854 28306 19906
rect 28306 19854 28308 19906
rect 28252 19852 28308 19854
rect 30716 19964 30772 20020
rect 29484 19852 29540 19908
rect 28588 19234 28644 19236
rect 28588 19182 28590 19234
rect 28590 19182 28642 19234
rect 28642 19182 28644 19234
rect 28588 19180 28644 19182
rect 29260 19234 29316 19236
rect 29260 19182 29262 19234
rect 29262 19182 29314 19234
rect 29314 19182 29316 19234
rect 29260 19180 29316 19182
rect 28364 18956 28420 19012
rect 30156 19180 30212 19236
rect 29372 18620 29428 18676
rect 27804 17948 27860 18004
rect 27244 16940 27300 16996
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 20860 40068 20916
rect 40012 19516 40068 19572
rect 37884 19292 37940 19348
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 30940 19010 30996 19012
rect 30940 18958 30942 19010
rect 30942 18958 30994 19010
rect 30994 18958 30996 19010
rect 30940 18956 30996 18958
rect 40012 18844 40068 18900
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 30268 16940 30324 16996
rect 27132 16882 27188 16884
rect 27132 16830 27134 16882
rect 27134 16830 27186 16882
rect 27186 16830 27188 16882
rect 27132 16828 27188 16830
rect 26348 16716 26404 16772
rect 26124 16658 26180 16660
rect 26124 16606 26126 16658
rect 26126 16606 26178 16658
rect 26178 16606 26180 16658
rect 26124 16604 26180 16606
rect 26348 16156 26404 16212
rect 27468 16716 27524 16772
rect 27804 16770 27860 16772
rect 27804 16718 27806 16770
rect 27806 16718 27858 16770
rect 27858 16718 27860 16770
rect 27804 16716 27860 16718
rect 26908 16492 26964 16548
rect 28476 16882 28532 16884
rect 28476 16830 28478 16882
rect 28478 16830 28530 16882
rect 28530 16830 28532 16882
rect 28476 16828 28532 16830
rect 37660 16882 37716 16884
rect 37660 16830 37662 16882
rect 37662 16830 37714 16882
rect 37714 16830 37716 16882
rect 37660 16828 37716 16830
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 39900 16156 39956 16212
rect 28028 16044 28084 16100
rect 37660 16098 37716 16100
rect 37660 16046 37662 16098
rect 37662 16046 37714 16098
rect 37714 16046 37716 16098
rect 37660 16044 37716 16046
rect 40012 15484 40068 15540
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 23548 5180 23604 5236
rect 20748 4114 20804 4116
rect 20748 4062 20750 4114
rect 20750 4062 20802 4114
rect 20802 4062 20804 4114
rect 20748 4060 20804 4062
rect 22876 3612 22932 3668
rect 20188 3388 20244 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21756 3388 21812 3444
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 24780 5234 24836 5236
rect 24780 5182 24782 5234
rect 24782 5182 24834 5234
rect 24834 5182 24836 5234
rect 24780 5180 24836 5182
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 25554 38556 25564 38612
rect 25620 38556 26796 38612
rect 26852 38556 26862 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 24882 38220 24892 38276
rect 24948 38220 26124 38276
rect 26180 38220 26190 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 21522 37436 21532 37492
rect 21588 37436 22764 37492
rect 22820 37436 22830 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 15474 36652 15484 36708
rect 15540 36652 16716 36708
rect 16772 36652 16782 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19506 28476 19516 28532
rect 19572 28476 20972 28532
rect 21028 28476 21038 28532
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 22530 28028 22540 28084
rect 22596 28028 23548 28084
rect 23604 28028 23614 28084
rect 17602 27804 17612 27860
rect 17668 27804 18172 27860
rect 18228 27804 19124 27860
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 19068 27524 19124 27804
rect 19058 27468 19068 27524
rect 19124 27468 19134 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 24546 27132 24556 27188
rect 24612 27132 25900 27188
rect 25956 27132 25966 27188
rect 4274 27020 4284 27076
rect 4340 27020 11788 27076
rect 11844 27020 11854 27076
rect 19506 27020 19516 27076
rect 19572 27020 20356 27076
rect 13346 26908 13356 26964
rect 13412 26908 14252 26964
rect 14308 26908 14318 26964
rect 17378 26908 17388 26964
rect 17444 26908 18844 26964
rect 18900 26908 19964 26964
rect 20020 26908 20030 26964
rect 20300 26852 20356 27020
rect 22418 26908 22428 26964
rect 22484 26908 23660 26964
rect 23716 26908 23726 26964
rect 20290 26796 20300 26852
rect 20356 26796 20366 26852
rect 20850 26796 20860 26852
rect 20916 26796 22204 26852
rect 22260 26796 22270 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 20178 26460 20188 26516
rect 20244 26460 21420 26516
rect 21476 26460 21486 26516
rect 23874 26460 23884 26516
rect 23940 26460 25788 26516
rect 25844 26460 25854 26516
rect 19618 26348 19628 26404
rect 19684 26348 20524 26404
rect 20580 26348 20748 26404
rect 20804 26348 20814 26404
rect 0 26292 800 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 14354 26236 14364 26292
rect 14420 26236 16156 26292
rect 16212 26236 16222 26292
rect 22530 26236 22540 26292
rect 22596 26236 23660 26292
rect 23716 26236 23726 26292
rect 23986 26236 23996 26292
rect 24052 26236 24444 26292
rect 24500 26236 24510 26292
rect 0 26208 800 26236
rect 15810 26124 15820 26180
rect 15876 26124 17388 26180
rect 17444 26124 17454 26180
rect 22978 26124 22988 26180
rect 23044 26124 23772 26180
rect 23828 26124 23838 26180
rect 23090 26012 23100 26068
rect 23156 26012 23660 26068
rect 23716 26012 23726 26068
rect 14914 25900 14924 25956
rect 14980 25900 15932 25956
rect 15988 25900 22652 25956
rect 22708 25900 23996 25956
rect 24052 25900 24062 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 22306 25564 22316 25620
rect 22372 25564 23324 25620
rect 23380 25564 23390 25620
rect 11778 25452 11788 25508
rect 11844 25452 14700 25508
rect 14756 25452 14766 25508
rect 16370 25452 16380 25508
rect 16436 25452 17500 25508
rect 17556 25452 17566 25508
rect 17938 25452 17948 25508
rect 18004 25452 18956 25508
rect 19012 25452 19022 25508
rect 16258 25340 16268 25396
rect 16324 25340 20076 25396
rect 20132 25340 20300 25396
rect 20356 25340 22428 25396
rect 22484 25340 22494 25396
rect 15362 25228 15372 25284
rect 15428 25228 16380 25284
rect 16436 25228 16446 25284
rect 17266 25228 17276 25284
rect 17332 25228 19180 25284
rect 19236 25228 22316 25284
rect 22372 25228 22382 25284
rect 22530 25228 22540 25284
rect 22596 25228 23436 25284
rect 23492 25228 23502 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 18946 24892 18956 24948
rect 19012 24892 20524 24948
rect 20580 24892 20590 24948
rect 12674 24668 12684 24724
rect 12740 24668 14588 24724
rect 14644 24668 15148 24724
rect 15204 24668 15708 24724
rect 15764 24668 15774 24724
rect 16482 24668 16492 24724
rect 16548 24668 18732 24724
rect 18788 24668 19180 24724
rect 19236 24668 19246 24724
rect 20738 24668 20748 24724
rect 20804 24668 22316 24724
rect 22372 24668 22382 24724
rect 28242 24668 28252 24724
rect 28308 24668 29484 24724
rect 29540 24668 37660 24724
rect 37716 24668 37726 24724
rect 18498 24444 18508 24500
rect 18564 24444 18956 24500
rect 19012 24444 19022 24500
rect 19618 24332 19628 24388
rect 19684 24332 20188 24388
rect 20244 24332 25900 24388
rect 25956 24332 25966 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 25890 23660 25900 23716
rect 25956 23660 27468 23716
rect 27524 23660 27534 23716
rect 41200 23604 42000 23632
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 22642 23436 22652 23492
rect 22708 23436 24556 23492
rect 24612 23436 24622 23492
rect 12002 23324 12012 23380
rect 12068 23324 20300 23380
rect 20356 23324 20860 23380
rect 20916 23324 20926 23380
rect 30034 23324 30044 23380
rect 30100 23324 37660 23380
rect 37716 23324 37726 23380
rect 15250 23212 15260 23268
rect 15316 23212 17388 23268
rect 17444 23212 17454 23268
rect 18610 23212 18620 23268
rect 18676 23212 18956 23268
rect 19012 23212 19022 23268
rect 27346 23212 27356 23268
rect 27412 23212 28364 23268
rect 28420 23212 28430 23268
rect 17714 23100 17724 23156
rect 17780 23100 19068 23156
rect 19124 23100 19134 23156
rect 19954 23100 19964 23156
rect 20020 23100 20636 23156
rect 20692 23100 20702 23156
rect 26852 23100 37660 23156
rect 37716 23100 37726 23156
rect 18722 22988 18732 23044
rect 18788 22988 19628 23044
rect 19684 22988 19694 23044
rect 26852 22932 26908 23100
rect 41200 22932 42000 22960
rect 24434 22876 24444 22932
rect 24500 22876 24668 22932
rect 24724 22876 26908 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14130 22540 14140 22596
rect 14196 22540 14924 22596
rect 14980 22540 14990 22596
rect 18610 22540 18620 22596
rect 18676 22540 19572 22596
rect 14924 22484 14980 22540
rect 19516 22484 19572 22540
rect 14924 22428 16380 22484
rect 16436 22428 18172 22484
rect 18228 22428 18956 22484
rect 19012 22428 19022 22484
rect 19506 22428 19516 22484
rect 19572 22428 21308 22484
rect 21364 22428 21374 22484
rect 26852 22428 27020 22484
rect 27076 22428 29596 22484
rect 29652 22428 29662 22484
rect 26852 22372 26908 22428
rect 14130 22316 14140 22372
rect 14196 22316 15372 22372
rect 15428 22316 16156 22372
rect 16212 22316 17388 22372
rect 17444 22316 18508 22372
rect 18564 22316 18574 22372
rect 19058 22316 19068 22372
rect 19124 22316 19292 22372
rect 19348 22316 26908 22372
rect 27458 22316 27468 22372
rect 27524 22316 30044 22372
rect 30100 22316 37660 22372
rect 37716 22316 37726 22372
rect 41200 22260 42000 22288
rect 20626 22204 20636 22260
rect 20692 22204 21644 22260
rect 21700 22204 21710 22260
rect 22642 22204 22652 22260
rect 22708 22204 24780 22260
rect 24836 22204 27356 22260
rect 27412 22204 29036 22260
rect 29092 22204 29102 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 12114 22092 12124 22148
rect 12180 22092 13916 22148
rect 13972 22092 14924 22148
rect 14980 22092 14990 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 17826 21868 17836 21924
rect 17892 21868 18284 21924
rect 18340 21868 19180 21924
rect 19236 21868 19246 21924
rect 17490 21644 17500 21700
rect 17556 21644 17948 21700
rect 18004 21644 20076 21700
rect 20132 21644 20142 21700
rect 26562 21532 26572 21588
rect 26628 21532 27132 21588
rect 27188 21532 27198 21588
rect 4162 21420 4172 21476
rect 4228 21420 16828 21476
rect 16884 21420 19404 21476
rect 19460 21420 19470 21476
rect 20066 21420 20076 21476
rect 20132 21420 23324 21476
rect 23380 21420 23390 21476
rect 23874 21196 23884 21252
rect 23940 21196 25228 21252
rect 25284 21196 25294 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 22642 20972 22652 21028
rect 22708 20972 23212 21028
rect 23268 20972 23278 21028
rect 41200 20916 42000 20944
rect 15138 20860 15148 20916
rect 15204 20860 17948 20916
rect 18004 20860 18014 20916
rect 22754 20860 22764 20916
rect 22820 20860 25340 20916
rect 25396 20860 26572 20916
rect 26628 20860 27468 20916
rect 27524 20860 27534 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 22642 20748 22652 20804
rect 22708 20748 24220 20804
rect 24276 20748 24286 20804
rect 15474 20636 15484 20692
rect 15540 20636 21532 20692
rect 21588 20636 22316 20692
rect 22372 20636 22382 20692
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 17826 20300 17836 20356
rect 17892 20300 19404 20356
rect 19460 20300 19470 20356
rect 19404 20244 19460 20300
rect 18722 20188 18732 20244
rect 18788 20188 19068 20244
rect 19124 20188 19134 20244
rect 19404 20188 21420 20244
rect 21476 20188 21486 20244
rect 22978 20076 22988 20132
rect 23044 20076 23772 20132
rect 23828 20076 28588 20132
rect 28644 20076 28654 20132
rect 14130 19964 14140 20020
rect 14196 19964 15260 20020
rect 15316 19964 15326 20020
rect 19170 19964 19180 20020
rect 19236 19964 20412 20020
rect 20468 19964 21308 20020
rect 21364 19964 21374 20020
rect 30706 19964 30716 20020
rect 30772 19964 37660 20020
rect 37716 19964 37726 20020
rect 12002 19852 12012 19908
rect 12068 19852 14476 19908
rect 14532 19852 14542 19908
rect 28242 19852 28252 19908
rect 28308 19852 29484 19908
rect 29540 19852 29550 19908
rect 18722 19740 18732 19796
rect 18788 19740 19740 19796
rect 19796 19740 19806 19796
rect 15586 19628 15596 19684
rect 15652 19628 16044 19684
rect 16100 19628 18620 19684
rect 18676 19628 20300 19684
rect 20356 19628 21644 19684
rect 21700 19628 21710 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 14578 19404 14588 19460
rect 14644 19404 15932 19460
rect 15988 19404 21756 19460
rect 21812 19404 21822 19460
rect 25778 19292 25788 19348
rect 25844 19292 37884 19348
rect 37940 19292 37950 19348
rect 28578 19180 28588 19236
rect 28644 19180 29260 19236
rect 29316 19180 29326 19236
rect 30146 19180 30156 19236
rect 30212 19180 37660 19236
rect 37716 19180 37726 19236
rect 16482 19068 16492 19124
rect 16548 19068 17052 19124
rect 17108 19068 17388 19124
rect 17444 19068 17612 19124
rect 17668 19068 17678 19124
rect 17938 19068 17948 19124
rect 18004 19068 26180 19124
rect 26124 19012 26180 19068
rect 11330 18956 11340 19012
rect 11396 18956 13804 19012
rect 13860 18956 14700 19012
rect 14756 18956 15372 19012
rect 15428 18956 17500 19012
rect 17556 18956 17566 19012
rect 17826 18956 17836 19012
rect 17892 18956 22316 19012
rect 22372 18956 23100 19012
rect 23156 18956 23166 19012
rect 26114 18956 26124 19012
rect 26180 18956 26908 19012
rect 26964 18956 26974 19012
rect 27122 18956 27132 19012
rect 27188 18956 27198 19012
rect 28354 18956 28364 19012
rect 28420 18956 30940 19012
rect 30996 18956 31006 19012
rect 17836 18900 17892 18956
rect 14018 18844 14028 18900
rect 14084 18844 14588 18900
rect 14644 18844 17892 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 27132 18788 27188 18956
rect 41200 18900 42000 18928
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 41200 18816 42000 18844
rect 14690 18732 14700 18788
rect 14756 18732 17724 18788
rect 17780 18732 17948 18788
rect 18004 18732 18014 18788
rect 26338 18732 26348 18788
rect 26404 18732 27188 18788
rect 15250 18620 15260 18676
rect 15316 18620 16716 18676
rect 16772 18620 18508 18676
rect 18564 18620 18574 18676
rect 26450 18620 26460 18676
rect 26516 18620 29372 18676
rect 29428 18620 29438 18676
rect 14466 18508 14476 18564
rect 14532 18508 15708 18564
rect 15764 18508 15774 18564
rect 4274 18396 4284 18452
rect 4340 18396 10668 18452
rect 10724 18396 14252 18452
rect 14308 18396 14318 18452
rect 17938 18396 17948 18452
rect 18004 18396 18620 18452
rect 18676 18396 19404 18452
rect 19460 18396 19470 18452
rect 20850 18396 20860 18452
rect 20916 18396 23324 18452
rect 23380 18396 23390 18452
rect 12338 18284 12348 18340
rect 12404 18284 14140 18340
rect 14196 18284 14206 18340
rect 16818 18284 16828 18340
rect 16884 18284 18172 18340
rect 18228 18284 18508 18340
rect 18564 18284 19292 18340
rect 19348 18284 19358 18340
rect 0 18228 800 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 0 18144 800 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 25666 17948 25676 18004
rect 25732 17948 27804 18004
rect 27860 17948 27870 18004
rect 18050 17836 18060 17892
rect 18116 17836 19068 17892
rect 19124 17836 19134 17892
rect 19618 17836 19628 17892
rect 19684 17836 22204 17892
rect 22260 17836 22270 17892
rect 16370 17612 16380 17668
rect 16436 17612 17724 17668
rect 17780 17612 17790 17668
rect 18946 17612 18956 17668
rect 19012 17612 19022 17668
rect 21858 17612 21868 17668
rect 21924 17612 22876 17668
rect 22932 17612 22942 17668
rect 18956 17444 19012 17612
rect 19618 17500 19628 17556
rect 19684 17500 20860 17556
rect 20916 17500 20926 17556
rect 16818 17388 16828 17444
rect 16884 17388 18396 17444
rect 18452 17388 19684 17444
rect 19628 17332 19684 17388
rect 19618 17276 19628 17332
rect 19684 17276 19694 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 18722 17164 18732 17220
rect 18788 17164 19684 17220
rect 22642 17164 22652 17220
rect 22708 17164 24556 17220
rect 24612 17164 24622 17220
rect 19628 17108 19684 17164
rect 19628 17052 20132 17108
rect 21410 17052 21420 17108
rect 21476 17052 25788 17108
rect 25844 17052 26908 17108
rect 26964 17052 26974 17108
rect 20076 16996 20132 17052
rect 14242 16940 14252 16996
rect 14308 16940 15036 16996
rect 15092 16940 15102 16996
rect 17154 16940 17164 16996
rect 17220 16940 19124 16996
rect 20076 16940 22764 16996
rect 22820 16940 26460 16996
rect 26516 16940 27244 16996
rect 27300 16940 27310 16996
rect 28252 16940 30268 16996
rect 30324 16940 30334 16996
rect 19068 16884 19124 16940
rect 28252 16884 28308 16940
rect 4274 16828 4284 16884
rect 4340 16828 12460 16884
rect 12516 16828 12526 16884
rect 15362 16828 15372 16884
rect 15428 16828 15708 16884
rect 15764 16828 17388 16884
rect 17444 16828 17454 16884
rect 18050 16828 18060 16884
rect 18116 16828 18732 16884
rect 18788 16828 18798 16884
rect 19068 16828 19740 16884
rect 19796 16828 22428 16884
rect 22484 16828 23212 16884
rect 23268 16828 23278 16884
rect 24546 16828 24556 16884
rect 24612 16828 27132 16884
rect 27188 16828 28308 16884
rect 28466 16828 28476 16884
rect 28532 16828 37660 16884
rect 37716 16828 37726 16884
rect 15474 16716 15484 16772
rect 15540 16716 16268 16772
rect 16324 16716 16604 16772
rect 16660 16716 17276 16772
rect 17332 16716 17342 16772
rect 26338 16716 26348 16772
rect 26404 16716 27468 16772
rect 27524 16716 27534 16772
rect 27794 16716 27804 16772
rect 27860 16716 27870 16772
rect 27804 16660 27860 16716
rect 14914 16604 14924 16660
rect 14980 16604 16492 16660
rect 16548 16604 16558 16660
rect 20066 16604 20076 16660
rect 20132 16604 21084 16660
rect 21140 16604 21150 16660
rect 26114 16604 26124 16660
rect 26180 16604 27860 16660
rect 15810 16492 15820 16548
rect 15876 16492 17612 16548
rect 17668 16492 18284 16548
rect 18340 16492 18350 16548
rect 26898 16492 26908 16548
rect 26964 16492 27002 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16212 800 16240
rect 41200 16212 42000 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 20402 16156 20412 16212
rect 20468 16156 23884 16212
rect 23940 16156 26348 16212
rect 26404 16156 26414 16212
rect 39890 16156 39900 16212
rect 39956 16156 42000 16212
rect 0 16128 800 16156
rect 41200 16128 42000 16156
rect 28018 16044 28028 16100
rect 28084 16044 37660 16100
rect 37716 16044 37726 16100
rect 12450 15932 12460 15988
rect 12516 15932 15596 15988
rect 15652 15932 15662 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 41200 15540 42000 15568
rect 18722 15484 18732 15540
rect 18788 15484 18798 15540
rect 40002 15484 40012 15540
rect 40068 15484 42000 15540
rect 18732 15204 18788 15484
rect 41200 15456 42000 15484
rect 14018 15148 14028 15204
rect 14084 15148 15708 15204
rect 15764 15148 15774 15204
rect 17602 15148 17612 15204
rect 17668 15148 20524 15204
rect 20580 15148 20590 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 18722 14588 18732 14644
rect 18788 14588 19628 14644
rect 19684 14588 19694 14644
rect 15586 14252 15596 14308
rect 15652 14252 17500 14308
rect 17556 14252 17566 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 17490 13692 17500 13748
rect 17556 13692 20748 13748
rect 20804 13692 20814 13748
rect 18498 13468 18508 13524
rect 18564 13468 19404 13524
rect 19460 13468 20300 13524
rect 20356 13468 20366 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 23538 5180 23548 5236
rect 23604 5180 24780 5236
rect 24836 5180 24846 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 19842 4060 19852 4116
rect 19908 4060 20748 4116
rect 20804 4060 20814 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 22866 3612 22876 3668
rect 22932 3612 25564 3668
rect 25620 3612 25630 3668
rect 20178 3388 20188 3444
rect 20244 3388 21756 3444
rect 21812 3388 21822 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 26908 17052 26964 17108
rect 26908 16492 26964 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 26908 17108 26964 17118
rect 26908 16548 26964 17052
rect 26908 16482 26964 16492
rect 35168 16492 35488 18004
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17584 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1698175906
transform 1 0 18256 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17136 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _106_
timestamp 1698175906
transform 1 0 14448 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26880 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 15120 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform 1 0 22176 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _112_
timestamp 1698175906
transform 1 0 27216 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _113_
timestamp 1698175906
transform -1 0 28336 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _114_
timestamp 1698175906
transform 1 0 17920 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform 1 0 18816 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform -1 0 18816 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _119_
timestamp 1698175906
transform -1 0 18144 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _120_
timestamp 1698175906
transform -1 0 17248 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform -1 0 20944 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_
timestamp 1698175906
transform -1 0 19824 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19600 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _124_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 -1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24976 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _128_
timestamp 1698175906
transform -1 0 22848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 23184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 23296 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _134_
timestamp 1698175906
transform -1 0 24080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24080 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform -1 0 23632 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform 1 0 20384 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15680 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14448 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _140_
timestamp 1698175906
transform -1 0 16576 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _141_
timestamp 1698175906
transform -1 0 16688 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1698175906
transform -1 0 18368 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform -1 0 15904 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 16240 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _145_
timestamp 1698175906
transform -1 0 15120 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _146_
timestamp 1698175906
transform -1 0 15008 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _148_
timestamp 1698175906
transform 1 0 14784 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _149_
timestamp 1698175906
transform 1 0 18032 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 18816
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13888 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _152_
timestamp 1698175906
transform 1 0 12208 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform 1 0 22176 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _154_
timestamp 1698175906
transform 1 0 17360 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _155_
timestamp 1698175906
transform -1 0 17920 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _156_
timestamp 1698175906
transform -1 0 15344 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _157_
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20384 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform -1 0 28560 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 27776 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _161_
timestamp 1698175906
transform -1 0 16688 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _162_
timestamp 1698175906
transform -1 0 16688 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1698175906
transform -1 0 14560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _164_
timestamp 1698175906
transform 1 0 19488 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1698175906
transform 1 0 20384 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _166_
timestamp 1698175906
transform -1 0 20384 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _167_
timestamp 1698175906
transform -1 0 19152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17136 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698175906
transform -1 0 18032 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _170_
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _171_
timestamp 1698175906
transform -1 0 28784 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform 1 0 20608 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _173_
timestamp 1698175906
transform 1 0 19712 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _174_
timestamp 1698175906
transform -1 0 18816 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _176_
timestamp 1698175906
transform 1 0 17248 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _177_
timestamp 1698175906
transform -1 0 16016 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16464 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _179_
timestamp 1698175906
transform 1 0 13888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform 1 0 24304 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform -1 0 22736 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform 1 0 23520 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _183_
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _184_
timestamp 1698175906
transform 1 0 22848 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _185_
timestamp 1698175906
transform 1 0 24080 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _186_
timestamp 1698175906
transform -1 0 28672 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _187_
timestamp 1698175906
transform 1 0 20720 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _188_
timestamp 1698175906
transform -1 0 27552 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform 1 0 30464 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26544 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _191_
timestamp 1698175906
transform 1 0 27888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25760 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _193_
timestamp 1698175906
transform -1 0 30464 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _194_
timestamp 1698175906
transform -1 0 29904 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _195_
timestamp 1698175906
transform -1 0 25536 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _196_
timestamp 1698175906
transform 1 0 14784 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698175906
transform 1 0 22176 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _198_
timestamp 1698175906
transform 1 0 22848 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _199_
timestamp 1698175906
transform 1 0 27552 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1698175906
transform -1 0 26320 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _201_
timestamp 1698175906
transform -1 0 22512 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _202_
timestamp 1698175906
transform 1 0 22064 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _203_
timestamp 1698175906
transform 1 0 22288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26992 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 21616 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 21616 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 11088 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 11200 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 11088 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform -1 0 13776 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 14896 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 26432 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 12432 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 17696 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 16016 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 26992 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 19152 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform -1 0 15568 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 22736 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 25536 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 27552 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 27328 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 22736 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 21504 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _232_
timestamp 1698175906
transform -1 0 23072 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _233_
timestamp 1698175906
transform 1 0 18816 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 14336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 14672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 15680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 17472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 20048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform -1 0 19152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 20720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 15568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 23184 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_312 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36288 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_328 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38080 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_336
timestamp 1698175906
transform 1 0 38976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_158
timestamp 1698175906
transform 1 0 19040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_162
timestamp 1698175906
transform 1 0 19488 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_189
timestamp 1698175906
transform 1 0 22512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_205
timestamp 1698175906
transform 1 0 24304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698175906
transform 1 0 22960 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_197
timestamp 1698175906
transform 1 0 23408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_225
timestamp 1698175906
transform 1 0 26544 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_171
timestamp 1698175906
transform 1 0 20496 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_175
timestamp 1698175906
transform 1 0 20944 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_111
timestamp 1698175906
transform 1 0 13776 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_116
timestamp 1698175906
transform 1 0 14336 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_124
timestamp 1698175906
transform 1 0 15232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_126
timestamp 1698175906
transform 1 0 15456 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_129
timestamp 1698175906
transform 1 0 15792 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_137
timestamp 1698175906
transform 1 0 16688 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_141
timestamp 1698175906
transform 1 0 17136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_143
timestamp 1698175906
transform 1 0 17360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_96
timestamp 1698175906
transform 1 0 12096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_135
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_176
timestamp 1698175906
transform 1 0 21056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_180
timestamp 1698175906
transform 1 0 21504 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_241
timestamp 1698175906
transform 1 0 28336 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_273
timestamp 1698175906
transform 1 0 31920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_131
timestamp 1698175906
transform 1 0 16016 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_141
timestamp 1698175906
transform 1 0 17136 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_153
timestamp 1698175906
transform 1 0 18480 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_169
timestamp 1698175906
transform 1 0 20272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_203
timestamp 1698175906
transform 1 0 24080 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_211
timestamp 1698175906
transform 1 0 24976 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_215
timestamp 1698175906
transform 1 0 25424 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_128
timestamp 1698175906
transform 1 0 15680 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_132
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_156
timestamp 1698175906
transform 1 0 18816 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_160
timestamp 1698175906
transform 1 0 19264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_168
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_172
timestamp 1698175906
transform 1 0 20608 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_181
timestamp 1698175906
transform 1 0 21616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_216
timestamp 1698175906
transform 1 0 25536 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_244
timestamp 1698175906
transform 1 0 28672 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698175906
transform 1 0 10864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_93
timestamp 1698175906
transform 1 0 11760 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_136
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_138
timestamp 1698175906
transform 1 0 16800 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_165
timestamp 1698175906
transform 1 0 19824 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_179
timestamp 1698175906
transform 1 0 21392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_209
timestamp 1698175906
transform 1 0 24752 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_111
timestamp 1698175906
transform 1 0 13776 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_122
timestamp 1698175906
transform 1 0 15008 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_130
timestamp 1698175906
transform 1 0 15904 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_175
timestamp 1698175906
transform 1 0 20944 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_183
timestamp 1698175906
transform 1 0 21840 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_201
timestamp 1698175906
transform 1 0 23856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698175906
transform 1 0 25536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_225
timestamp 1698175906
transform 1 0 26544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_227
timestamp 1698175906
transform 1 0 26768 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_233
timestamp 1698175906
transform 1 0 27440 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_263
timestamp 1698175906
transform 1 0 30800 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_113
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_133
timestamp 1698175906
transform 1 0 16240 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_189
timestamp 1698175906
transform 1 0 22512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_220
timestamp 1698175906
transform 1 0 25984 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_224
timestamp 1698175906
transform 1 0 26432 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_234
timestamp 1698175906
transform 1 0 27552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_236
timestamp 1698175906
transform 1 0 27776 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_265
timestamp 1698175906
transform 1 0 31024 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_297
timestamp 1698175906
transform 1 0 34608 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698175906
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_84
timestamp 1698175906
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_86
timestamp 1698175906
transform 1 0 10976 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_122
timestamp 1698175906
transform 1 0 15008 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_152
timestamp 1698175906
transform 1 0 18368 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_157
timestamp 1698175906
transform 1 0 18928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_202
timestamp 1698175906
transform 1 0 23968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_216
timestamp 1698175906
transform 1 0 25536 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_261
timestamp 1698175906
transform 1 0 30576 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_192
timestamp 1698175906
transform 1 0 22848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_194
timestamp 1698175906
transform 1 0 23072 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_117
timestamp 1698175906
transform 1 0 14448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_121
timestamp 1698175906
transform 1 0 14896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_123
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_130
timestamp 1698175906
transform 1 0 15904 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_157
timestamp 1698175906
transform 1 0 18928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_159
timestamp 1698175906
transform 1 0 19152 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_228
timestamp 1698175906
transform 1 0 26880 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_258
timestamp 1698175906
transform 1 0 30240 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 32032 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_117
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_119
timestamp 1698175906
transform 1 0 14672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_136
timestamp 1698175906
transform 1 0 16576 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_140
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_183
timestamp 1698175906
transform 1 0 21840 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_185
timestamp 1698175906
transform 1 0 22064 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_211
timestamp 1698175906
transform 1 0 24976 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_227
timestamp 1698175906
transform 1 0 26768 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_255
timestamp 1698175906
transform 1 0 29904 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_287
timestamp 1698175906
transform 1 0 33488 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_303
timestamp 1698175906
transform 1 0 35280 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_84
timestamp 1698175906
transform 1 0 10752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_86
timestamp 1698175906
transform 1 0 10976 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_128
timestamp 1698175906
transform 1 0 15680 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_156
timestamp 1698175906
transform 1 0 18816 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_176
timestamp 1698175906
transform 1 0 21056 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_180
timestamp 1698175906
transform 1 0 21504 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_228
timestamp 1698175906
transform 1 0 26880 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_258
timestamp 1698175906
transform 1 0 30240 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698175906
transform 1 0 32032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_118
timestamp 1698175906
transform 1 0 14560 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_150
timestamp 1698175906
transform 1 0 18144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_162
timestamp 1698175906
transform 1 0 19488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_170
timestamp 1698175906
transform 1 0 20384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698175906
transform 1 0 22288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_192
timestamp 1698175906
transform 1 0 22848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_224
timestamp 1698175906
transform 1 0 26432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_228
timestamp 1698175906
transform 1 0 26880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_230
timestamp 1698175906
transform 1 0 27104 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_236
timestamp 1698175906
transform 1 0 27776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_121
timestamp 1698175906
transform 1 0 14896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_125
timestamp 1698175906
transform 1 0 15344 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_133
timestamp 1698175906
transform 1 0 16240 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698175906
transform 1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_150
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_159
timestamp 1698175906
transform 1 0 19152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_167
timestamp 1698175906
transform 1 0 20048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_175
timestamp 1698175906
transform 1 0 20944 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_183
timestamp 1698175906
transform 1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_185
timestamp 1698175906
transform 1 0 22064 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_192
timestamp 1698175906
transform 1 0 22848 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_253
timestamp 1698175906
transform 1 0 29680 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_269
timestamp 1698175906
transform 1 0 31472 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_111
timestamp 1698175906
transform 1 0 13776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_115
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_125
timestamp 1698175906
transform 1 0 15344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_127
timestamp 1698175906
transform 1 0 15568 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_130
timestamp 1698175906
transform 1 0 15904 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_137
timestamp 1698175906
transform 1 0 16688 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_163
timestamp 1698175906
transform 1 0 19600 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_185
timestamp 1698175906
transform 1 0 22064 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_220
timestamp 1698175906
transform 1 0 25984 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_236
timestamp 1698175906
transform 1 0 27776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_96
timestamp 1698175906
transform 1 0 12096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_98
timestamp 1698175906
transform 1 0 12320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698175906
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_177
timestamp 1698175906
transform 1 0 21168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_181
timestamp 1698175906
transform 1 0 21616 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_189
timestamp 1698175906
transform 1 0 22512 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_191
timestamp 1698175906
transform 1 0 22736 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698175906
transform 1 0 14000 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_118
timestamp 1698175906
transform 1 0 14560 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_126
timestamp 1698175906
transform 1 0 15456 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_130
timestamp 1698175906
transform 1 0 15904 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_165
timestamp 1698175906
transform 1 0 19824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_169
timestamp 1698175906
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_189
timestamp 1698175906
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_191
timestamp 1698175906
transform 1 0 22736 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_221
timestamp 1698175906
transform 1 0 26096 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_237
timestamp 1698175906
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_149
timestamp 1698175906
transform 1 0 18032 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_194
timestamp 1698175906
transform 1 0 23072 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_203
timestamp 1698175906
transform 1 0 24080 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_123
timestamp 1698175906
transform 1 0 15120 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_153
timestamp 1698175906
transform 1 0 18480 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_169
timestamp 1698175906
transform 1 0 20272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 18592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 24864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 27888 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_256
timestamp 1698175906
transform 1 0 30016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_258
timestamp 1698175906
transform 1 0 30240 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_263
timestamp 1698175906
transform 1 0 30800 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698175906
transform 1 0 31696 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita1_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 30800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita1_26
timestamp 1698175906
transform -1 0 36288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 24192 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 19600 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 21616 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 24976 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 15568 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 21616 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 23632 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 30240 41200 30352 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 41200 15456 42000 15568 0 FreeSans 448 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 21504 41200 21616 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 15456 41200 15568 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 18200 14840 18200 14840 0 _000_
rlabel metal2 14168 14952 14168 14952 0 _001_
rlabel metal2 23800 27384 23800 27384 0 _002_
rlabel metal2 23688 25816 23688 25816 0 _003_
rlabel metal2 26544 16184 26544 16184 0 _004_
rlabel metal2 28504 18592 28504 18592 0 _005_
rlabel metal2 29512 19432 29512 19432 0 _006_
rlabel metal2 23744 22120 23744 22120 0 _007_
rlabel metal2 26040 16072 26040 16072 0 _008_
rlabel metal2 22512 17752 22512 17752 0 _009_
rlabel metal2 27888 21672 27888 21672 0 _010_
rlabel metal2 18256 26152 18256 26152 0 _011_
rlabel metal2 22568 23352 22568 23352 0 _012_
rlabel metal2 22568 15792 22568 15792 0 _013_
rlabel metal2 20328 24360 20328 24360 0 _014_
rlabel metal3 13048 22120 13048 22120 0 _015_
rlabel metal3 13272 19880 13272 19880 0 _016_
rlabel metal3 14672 16968 14672 16968 0 _017_
rlabel metal2 12488 18088 12488 18088 0 _018_
rlabel metal2 13944 25032 13944 25032 0 _019_
rlabel metal2 27440 24136 27440 24136 0 _020_
rlabel metal2 13384 26656 13384 26656 0 _021_
rlabel metal2 18648 14560 18648 14560 0 _022_
rlabel metal2 16968 27384 16968 27384 0 _023_
rlabel metal2 28504 22792 28504 22792 0 _024_
rlabel metal2 20440 26320 20440 26320 0 _025_
rlabel metal3 17640 24696 17640 24696 0 _026_
rlabel metal2 26152 18816 26152 18816 0 _027_
rlabel metal2 12376 18032 12376 18032 0 _028_
rlabel metal2 22680 25424 22680 25424 0 _029_
rlabel metal3 18424 23128 18424 23128 0 _030_
rlabel metal2 15176 25312 15176 25312 0 _031_
rlabel metal2 14056 25592 14056 25592 0 _032_
rlabel metal2 25928 24024 25928 24024 0 _033_
rlabel metal2 27832 23800 27832 23800 0 _034_
rlabel metal2 16296 25928 16296 25928 0 _035_
rlabel metal3 15288 26264 15288 26264 0 _036_
rlabel metal2 20216 16072 20216 16072 0 _037_
rlabel metal2 20552 15400 20552 15400 0 _038_
rlabel metal2 18424 24920 18424 24920 0 _039_
rlabel metal2 17864 26488 17864 26488 0 _040_
rlabel metal2 29288 22512 29288 22512 0 _041_
rlabel metal2 20664 25760 20664 25760 0 _042_
rlabel metal2 18536 15736 18536 15736 0 _043_
rlabel metal2 17696 16296 17696 16296 0 _044_
rlabel metal2 16072 15344 16072 15344 0 _045_
rlabel metal2 14056 14896 14056 14896 0 _046_
rlabel metal2 24472 26040 24472 26040 0 _047_
rlabel metal2 22456 26320 22456 26320 0 _048_
rlabel metal3 23408 26152 23408 26152 0 _049_
rlabel metal2 23856 22456 23856 22456 0 _050_
rlabel metal2 27384 17080 27384 17080 0 _051_
rlabel metal2 25816 16968 25816 16968 0 _052_
rlabel metal3 29680 18984 29680 18984 0 _053_
rlabel metal2 27944 19264 27944 19264 0 _054_
rlabel metal2 26488 18536 26488 18536 0 _055_
rlabel metal2 29848 19096 29848 19096 0 _056_
rlabel metal3 24584 21224 24584 21224 0 _057_
rlabel metal3 21952 20664 21952 20664 0 _058_
rlabel metal3 22960 21000 22960 21000 0 _059_
rlabel metal3 27832 16688 27832 16688 0 _060_
rlabel metal2 22120 19040 22120 19040 0 _061_
rlabel metal2 22344 17752 22344 17752 0 _062_
rlabel metal2 21448 20496 21448 20496 0 _063_
rlabel metal3 17640 17416 17640 17416 0 _064_
rlabel metal3 24640 16968 24640 16968 0 _065_
rlabel metal2 20440 19208 20440 19208 0 _066_
rlabel metal2 20216 22008 20216 22008 0 _067_
rlabel metal2 19320 22232 19320 22232 0 _068_
rlabel metal2 27384 20160 27384 20160 0 _069_
rlabel metal2 20328 18984 20328 18984 0 _070_
rlabel metal3 21560 24696 21560 24696 0 _071_
rlabel metal3 23744 22232 23744 22232 0 _072_
rlabel metal2 27944 22344 27944 22344 0 _073_
rlabel metal2 18648 22792 18648 22792 0 _074_
rlabel metal2 23408 26264 23408 26264 0 _075_
rlabel metal2 22232 17416 22232 17416 0 _076_
rlabel metal2 18200 18368 18200 18368 0 _077_
rlabel metal2 17640 16688 17640 16688 0 _078_
rlabel metal2 17080 18480 17080 18480 0 _079_
rlabel metal2 18648 24752 18648 24752 0 _080_
rlabel metal2 20552 25648 20552 25648 0 _081_
rlabel metal2 19376 25704 19376 25704 0 _082_
rlabel metal2 21784 22232 21784 22232 0 _083_
rlabel metal2 17640 15568 17640 15568 0 _084_
rlabel metal3 23464 20776 23464 20776 0 _085_
rlabel metal2 24584 22792 24584 22792 0 _086_
rlabel metal2 20888 17696 20888 17696 0 _087_
rlabel metal2 23464 22064 23464 22064 0 _088_
rlabel metal2 23016 17528 23016 17528 0 _089_
rlabel metal3 22848 16856 22848 16856 0 _090_
rlabel metal3 22176 16184 22176 16184 0 _091_
rlabel metal2 23968 17080 23968 17080 0 _092_
rlabel metal2 23464 16464 23464 16464 0 _093_
rlabel metal2 14280 22680 14280 22680 0 _094_
rlabel metal2 15736 21952 15736 21952 0 _095_
rlabel metal2 15960 19600 15960 19600 0 _096_
rlabel metal2 23072 22232 23072 22232 0 _097_
rlabel metal2 15232 21784 15232 21784 0 _098_
rlabel metal2 15400 16408 15400 16408 0 _099_
rlabel metal2 14840 19544 14840 19544 0 _100_
rlabel metal3 16072 16744 16072 16744 0 _101_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 23352 21112 23352 21112 0 clknet_0_clk
rlabel metal3 20832 26488 20832 26488 0 clknet_1_0__leaf_clk
rlabel metal2 22904 26264 22904 26264 0 clknet_1_1__leaf_clk
rlabel metal2 18200 22792 18200 22792 0 dut1.count\[0\]
rlabel metal3 17976 22344 17976 22344 0 dut1.count\[1\]
rlabel metal2 14560 20552 14560 20552 0 dut1.count\[2\]
rlabel metal2 16408 17696 16408 17696 0 dut1.count\[3\]
rlabel metal2 25368 19600 25368 19600 0 net1
rlabel metal2 30744 19544 30744 19544 0 net10
rlabel metal2 19096 27328 19096 27328 0 net11
rlabel metal2 30184 19152 30184 19152 0 net12
rlabel metal2 20720 3528 20720 3528 0 net13
rlabel metal2 24584 26824 24584 26824 0 net14
rlabel metal3 24864 26488 24864 26488 0 net15
rlabel metal2 16072 25984 16072 25984 0 net16
rlabel metal2 29512 24640 29512 24640 0 net17
rlabel metal2 11816 25816 11816 25816 0 net18
rlabel metal2 10696 18368 10696 18368 0 net19
rlabel metal2 30072 23184 30072 23184 0 net2
rlabel metal2 24696 22960 24696 22960 0 net20
rlabel metal3 20328 26936 20328 26936 0 net21
rlabel metal2 12488 16016 12488 16016 0 net22
rlabel metal2 30072 21896 30072 21896 0 net23
rlabel metal2 23800 6748 23800 6748 0 net24
rlabel metal2 30408 37912 30408 37912 0 net25
rlabel metal2 35672 2030 35672 2030 0 net26
rlabel metal2 28056 16464 28056 16464 0 net3
rlabel metal2 24584 5964 24584 5964 0 net4
rlabel metal3 23072 28056 23072 28056 0 net5
rlabel metal2 19712 4312 19712 4312 0 net6
rlabel metal2 20328 13552 20328 13552 0 net7
rlabel metal2 22456 27720 22456 27720 0 net8
rlabel metal3 33096 16856 33096 16856 0 net9
rlabel metal2 40040 21112 40040 21112 0 segm[10]
rlabel metal2 40040 23800 40040 23800 0 segm[11]
rlabel metal2 40040 15848 40040 15848 0 segm[12]
rlabel metal2 22904 2198 22904 2198 0 segm[13]
rlabel metal2 22232 39690 22232 39690 0 segm[1]
rlabel metal2 19544 2030 19544 2030 0 segm[2]
rlabel metal2 18872 2198 18872 2198 0 segm[3]
rlabel metal2 21560 39354 21560 39354 0 segm[4]
rlabel metal2 39928 16464 39928 16464 0 segm[6]
rlabel metal2 40040 19656 40040 19656 0 segm[7]
rlabel metal2 18872 39690 18872 39690 0 segm[8]
rlabel metal2 40040 19096 40040 19096 0 segm[9]
rlabel metal2 20216 2086 20216 2086 0 sel[0]
rlabel metal2 25592 39914 25592 39914 0 sel[10]
rlabel metal2 24920 39746 24920 39746 0 sel[11]
rlabel metal2 15512 38962 15512 38962 0 sel[1]
rlabel metal2 40040 24360 40040 24360 0 sel[2]
rlabel metal3 1358 26264 1358 26264 0 sel[3]
rlabel metal3 1358 18200 1358 18200 0 sel[4]
rlabel metal3 40642 22904 40642 22904 0 sel[5]
rlabel metal2 19544 39186 19544 39186 0 sel[6]
rlabel metal3 1358 16184 1358 16184 0 sel[7]
rlabel metal2 40040 22344 40040 22344 0 sel[8]
rlabel metal2 23576 2982 23576 2982 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
