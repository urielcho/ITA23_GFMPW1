magic
tech gf180mcuD
magscale 1 10
timestamp 1699642850
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 26798 37490 26850 37502
rect 26798 37426 26850 37438
rect 25778 37214 25790 37266
rect 25842 37214 25854 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 21422 28530 21474 28542
rect 21422 28466 21474 28478
rect 17838 28418 17890 28430
rect 17838 28354 17890 28366
rect 21310 28418 21362 28430
rect 21310 28354 21362 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 15262 28082 15314 28094
rect 15262 28018 15314 28030
rect 25342 28082 25394 28094
rect 25342 28018 25394 28030
rect 14702 27970 14754 27982
rect 14702 27906 14754 27918
rect 17950 27970 18002 27982
rect 17950 27906 18002 27918
rect 18734 27970 18786 27982
rect 23998 27970 24050 27982
rect 20850 27918 20862 27970
rect 20914 27918 20926 27970
rect 18734 27906 18786 27918
rect 23998 27906 24050 27918
rect 14478 27858 14530 27870
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 14242 27806 14254 27858
rect 14306 27806 14318 27858
rect 14478 27794 14530 27806
rect 14814 27858 14866 27870
rect 17614 27858 17666 27870
rect 17378 27806 17390 27858
rect 17442 27806 17454 27858
rect 14814 27794 14866 27806
rect 17614 27794 17666 27806
rect 17838 27858 17890 27870
rect 17838 27794 17890 27806
rect 18398 27858 18450 27870
rect 23774 27858 23826 27870
rect 20178 27806 20190 27858
rect 20242 27806 20254 27858
rect 18398 27794 18450 27806
rect 23774 27794 23826 27806
rect 24110 27858 24162 27870
rect 24110 27794 24162 27806
rect 25118 27858 25170 27870
rect 25118 27794 25170 27806
rect 25454 27858 25506 27870
rect 25454 27794 25506 27806
rect 16830 27746 16882 27758
rect 11330 27694 11342 27746
rect 11394 27694 11406 27746
rect 13458 27694 13470 27746
rect 13522 27694 13534 27746
rect 16830 27682 16882 27694
rect 17726 27746 17778 27758
rect 23438 27746 23490 27758
rect 22978 27694 22990 27746
rect 23042 27694 23054 27746
rect 17726 27682 17778 27694
rect 23438 27682 23490 27694
rect 1934 27634 1986 27646
rect 1934 27570 1986 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 27470 27298 27522 27310
rect 27470 27234 27522 27246
rect 1934 27186 1986 27198
rect 21646 27186 21698 27198
rect 40014 27186 40066 27198
rect 15362 27134 15374 27186
rect 15426 27134 15438 27186
rect 17490 27134 17502 27186
rect 17554 27134 17566 27186
rect 18610 27134 18622 27186
rect 18674 27134 18686 27186
rect 20738 27134 20750 27186
rect 20802 27134 20814 27186
rect 23762 27134 23774 27186
rect 23826 27134 23838 27186
rect 25890 27134 25902 27186
rect 25954 27134 25966 27186
rect 1934 27122 1986 27134
rect 21646 27122 21698 27134
rect 40014 27122 40066 27134
rect 14366 27074 14418 27086
rect 21534 27074 21586 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 14578 27022 14590 27074
rect 14642 27022 14654 27074
rect 17938 27022 17950 27074
rect 18002 27022 18014 27074
rect 21298 27022 21310 27074
rect 21362 27022 21374 27074
rect 14366 27010 14418 27022
rect 21534 27010 21586 27022
rect 21758 27074 21810 27086
rect 27134 27074 27186 27086
rect 21970 27022 21982 27074
rect 22034 27022 22046 27074
rect 22978 27022 22990 27074
rect 23042 27022 23054 27074
rect 21758 27010 21810 27022
rect 27134 27010 27186 27022
rect 27582 27074 27634 27086
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 27582 27010 27634 27022
rect 13918 26962 13970 26974
rect 13918 26898 13970 26910
rect 26798 26962 26850 26974
rect 26798 26898 26850 26910
rect 26910 26962 26962 26974
rect 26910 26898 26962 26910
rect 13694 26850 13746 26862
rect 13694 26786 13746 26798
rect 13806 26850 13858 26862
rect 13806 26786 13858 26798
rect 26350 26850 26402 26862
rect 26350 26786 26402 26798
rect 27470 26850 27522 26862
rect 27470 26786 27522 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 15150 26514 15202 26526
rect 15150 26450 15202 26462
rect 15822 26514 15874 26526
rect 15822 26450 15874 26462
rect 20974 26514 21026 26526
rect 24670 26514 24722 26526
rect 21970 26462 21982 26514
rect 22034 26462 22046 26514
rect 20974 26450 21026 26462
rect 24670 26450 24722 26462
rect 16046 26402 16098 26414
rect 18510 26402 18562 26414
rect 13906 26350 13918 26402
rect 13970 26350 13982 26402
rect 16482 26350 16494 26402
rect 16546 26350 16558 26402
rect 16046 26338 16098 26350
rect 18510 26338 18562 26350
rect 18846 26402 18898 26414
rect 18846 26338 18898 26350
rect 18958 26402 19010 26414
rect 18958 26338 19010 26350
rect 23662 26402 23714 26414
rect 26226 26350 26238 26402
rect 26290 26350 26302 26402
rect 23662 26338 23714 26350
rect 14926 26290 14978 26302
rect 14578 26238 14590 26290
rect 14642 26238 14654 26290
rect 14926 26226 14978 26238
rect 15262 26290 15314 26302
rect 15262 26226 15314 26238
rect 16158 26290 16210 26302
rect 16158 26226 16210 26238
rect 16830 26290 16882 26302
rect 19518 26290 19570 26302
rect 23550 26290 23602 26302
rect 17826 26238 17838 26290
rect 17890 26238 17902 26290
rect 19170 26238 19182 26290
rect 19234 26238 19246 26290
rect 21746 26238 21758 26290
rect 21810 26238 21822 26290
rect 16830 26226 16882 26238
rect 19518 26226 19570 26238
rect 23550 26226 23602 26238
rect 23886 26290 23938 26302
rect 25442 26238 25454 26290
rect 25506 26238 25518 26290
rect 23886 26226 23938 26238
rect 11778 26126 11790 26178
rect 11842 26126 11854 26178
rect 17602 26126 17614 26178
rect 17666 26126 17678 26178
rect 28354 26126 28366 26178
rect 28418 26126 28430 26178
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 17614 25730 17666 25742
rect 17614 25666 17666 25678
rect 13582 25618 13634 25630
rect 13582 25554 13634 25566
rect 14926 25618 14978 25630
rect 14926 25554 14978 25566
rect 19294 25618 19346 25630
rect 26238 25618 26290 25630
rect 22866 25566 22878 25618
rect 22930 25566 22942 25618
rect 24994 25566 25006 25618
rect 25058 25566 25070 25618
rect 19294 25554 19346 25566
rect 26238 25554 26290 25566
rect 40014 25618 40066 25630
rect 40014 25554 40066 25566
rect 13470 25506 13522 25518
rect 13470 25442 13522 25454
rect 14142 25506 14194 25518
rect 14142 25442 14194 25454
rect 16158 25506 16210 25518
rect 27022 25506 27074 25518
rect 18162 25454 18174 25506
rect 18226 25454 18238 25506
rect 19954 25454 19966 25506
rect 20018 25454 20030 25506
rect 25666 25454 25678 25506
rect 25730 25454 25742 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 16158 25442 16210 25454
rect 27022 25442 27074 25454
rect 16382 25394 16434 25406
rect 16382 25330 16434 25342
rect 16494 25394 16546 25406
rect 16494 25330 16546 25342
rect 17726 25394 17778 25406
rect 17726 25330 17778 25342
rect 17950 25394 18002 25406
rect 17950 25330 18002 25342
rect 19182 25394 19234 25406
rect 19182 25330 19234 25342
rect 19406 25394 19458 25406
rect 19406 25330 19458 25342
rect 27134 25394 27186 25406
rect 27134 25330 27186 25342
rect 13694 25282 13746 25294
rect 13694 25218 13746 25230
rect 16942 25282 16994 25294
rect 16942 25218 16994 25230
rect 17390 25282 17442 25294
rect 27358 25282 27410 25294
rect 19730 25230 19742 25282
rect 19794 25230 19806 25282
rect 17390 25218 17442 25230
rect 27358 25218 27410 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 18622 24946 18674 24958
rect 18274 24894 18286 24946
rect 18338 24894 18350 24946
rect 18622 24882 18674 24894
rect 25454 24946 25506 24958
rect 25454 24882 25506 24894
rect 22978 24782 22990 24834
rect 23042 24782 23054 24834
rect 19506 24670 19518 24722
rect 19570 24670 19582 24722
rect 25778 24670 25790 24722
rect 25842 24670 25854 24722
rect 26562 24558 26574 24610
rect 26626 24558 26638 24610
rect 28690 24558 28702 24610
rect 28754 24558 28766 24610
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 23662 24162 23714 24174
rect 23662 24098 23714 24110
rect 26462 24162 26514 24174
rect 26462 24098 26514 24110
rect 1934 24050 1986 24062
rect 17614 24050 17666 24062
rect 25342 24050 25394 24062
rect 16370 23998 16382 24050
rect 16434 23998 16446 24050
rect 21858 23998 21870 24050
rect 21922 23998 21934 24050
rect 24770 23998 24782 24050
rect 24834 23998 24846 24050
rect 1934 23986 1986 23998
rect 17614 23986 17666 23998
rect 25342 23986 25394 23998
rect 16830 23938 16882 23950
rect 21422 23938 21474 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 13570 23886 13582 23938
rect 13634 23886 13646 23938
rect 20626 23886 20638 23938
rect 20690 23886 20702 23938
rect 16830 23874 16882 23886
rect 21422 23874 21474 23886
rect 22318 23938 22370 23950
rect 22318 23874 22370 23886
rect 24334 23938 24386 23950
rect 24334 23874 24386 23886
rect 26574 23938 26626 23950
rect 26574 23874 26626 23886
rect 23214 23826 23266 23838
rect 14242 23774 14254 23826
rect 14306 23774 14318 23826
rect 20290 23774 20302 23826
rect 20354 23774 20366 23826
rect 22866 23774 22878 23826
rect 22930 23774 22942 23826
rect 23214 23762 23266 23774
rect 23774 23826 23826 23838
rect 23774 23762 23826 23774
rect 21310 23714 21362 23726
rect 17154 23662 17166 23714
rect 17218 23662 17230 23714
rect 20626 23662 20638 23714
rect 20690 23662 20702 23714
rect 21310 23650 21362 23662
rect 23662 23714 23714 23726
rect 23662 23650 23714 23662
rect 26462 23714 26514 23726
rect 26462 23650 26514 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 14366 23378 14418 23390
rect 14366 23314 14418 23326
rect 17726 23378 17778 23390
rect 17726 23314 17778 23326
rect 18958 23378 19010 23390
rect 18958 23314 19010 23326
rect 21870 23378 21922 23390
rect 21870 23314 21922 23326
rect 24222 23378 24274 23390
rect 24222 23314 24274 23326
rect 22990 23266 23042 23278
rect 18610 23214 18622 23266
rect 18674 23214 18686 23266
rect 22990 23202 23042 23214
rect 14478 23154 14530 23166
rect 13682 23102 13694 23154
rect 13746 23102 13758 23154
rect 14478 23090 14530 23102
rect 15374 23154 15426 23166
rect 15374 23090 15426 23102
rect 20862 23154 20914 23166
rect 22766 23154 22818 23166
rect 21746 23102 21758 23154
rect 21810 23102 21822 23154
rect 20862 23090 20914 23102
rect 22766 23090 22818 23102
rect 23662 23154 23714 23166
rect 24434 23102 24446 23154
rect 24498 23102 24510 23154
rect 28242 23102 28254 23154
rect 28306 23102 28318 23154
rect 23662 23090 23714 23102
rect 15710 23042 15762 23054
rect 10882 22990 10894 23042
rect 10946 22990 10958 23042
rect 13010 22990 13022 23042
rect 13074 22990 13086 23042
rect 15710 22978 15762 22990
rect 18286 23042 18338 23054
rect 19966 23042 20018 23054
rect 19618 22990 19630 23042
rect 19682 22990 19694 23042
rect 20402 22990 20414 23042
rect 20466 22990 20478 23042
rect 21522 22990 21534 23042
rect 21586 22990 21598 23042
rect 25442 22990 25454 23042
rect 25506 22990 25518 23042
rect 27570 22990 27582 23042
rect 27634 22990 27646 23042
rect 18286 22978 18338 22990
rect 19966 22978 20018 22990
rect 14366 22930 14418 22942
rect 14366 22866 14418 22878
rect 15150 22930 15202 22942
rect 15150 22866 15202 22878
rect 15262 22930 15314 22942
rect 15262 22866 15314 22878
rect 15934 22930 15986 22942
rect 15934 22866 15986 22878
rect 22430 22930 22482 22942
rect 22430 22866 22482 22878
rect 23326 22930 23378 22942
rect 23326 22866 23378 22878
rect 23438 22930 23490 22942
rect 23438 22866 23490 22878
rect 23774 22930 23826 22942
rect 23774 22866 23826 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 17278 22594 17330 22606
rect 17278 22530 17330 22542
rect 17950 22594 18002 22606
rect 17950 22530 18002 22542
rect 25230 22594 25282 22606
rect 25230 22530 25282 22542
rect 26350 22594 26402 22606
rect 26350 22530 26402 22542
rect 1934 22482 1986 22494
rect 1934 22418 1986 22430
rect 14030 22482 14082 22494
rect 19282 22430 19294 22482
rect 19346 22430 19358 22482
rect 14030 22418 14082 22430
rect 17166 22370 17218 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 17166 22306 17218 22318
rect 17726 22370 17778 22382
rect 17726 22306 17778 22318
rect 18286 22370 18338 22382
rect 18286 22306 18338 22318
rect 20190 22370 20242 22382
rect 20190 22306 20242 22318
rect 20750 22370 20802 22382
rect 25118 22370 25170 22382
rect 22866 22318 22878 22370
rect 22930 22318 22942 22370
rect 24770 22318 24782 22370
rect 24834 22318 24846 22370
rect 20750 22306 20802 22318
rect 25118 22306 25170 22318
rect 25678 22370 25730 22382
rect 25678 22306 25730 22318
rect 18510 22258 18562 22270
rect 24894 22258 24946 22270
rect 22082 22206 22094 22258
rect 22146 22206 22158 22258
rect 23090 22206 23102 22258
rect 23154 22206 23166 22258
rect 18510 22194 18562 22206
rect 24894 22194 24946 22206
rect 26238 22258 26290 22270
rect 26238 22194 26290 22206
rect 17614 22146 17666 22158
rect 17614 22082 17666 22094
rect 18846 22146 18898 22158
rect 18846 22082 18898 22094
rect 19854 22146 19906 22158
rect 19854 22082 19906 22094
rect 25230 22146 25282 22158
rect 25230 22082 25282 22094
rect 25790 22146 25842 22158
rect 25790 22082 25842 22094
rect 26014 22146 26066 22158
rect 26014 22082 26066 22094
rect 26350 22146 26402 22158
rect 26350 22082 26402 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14030 21810 14082 21822
rect 14030 21746 14082 21758
rect 14702 21810 14754 21822
rect 14702 21746 14754 21758
rect 19070 21698 19122 21710
rect 40238 21698 40290 21710
rect 12786 21646 12798 21698
rect 12850 21646 12862 21698
rect 15250 21646 15262 21698
rect 15314 21646 15326 21698
rect 15810 21646 15822 21698
rect 15874 21646 15886 21698
rect 18162 21646 18174 21698
rect 18226 21646 18238 21698
rect 18498 21646 18510 21698
rect 18562 21646 18574 21698
rect 25554 21646 25566 21698
rect 25618 21646 25630 21698
rect 19070 21634 19122 21646
rect 40238 21634 40290 21646
rect 15486 21586 15538 21598
rect 13570 21534 13582 21586
rect 13634 21534 13646 21586
rect 14914 21534 14926 21586
rect 14978 21534 14990 21586
rect 15486 21522 15538 21534
rect 16158 21586 16210 21598
rect 16482 21534 16494 21586
rect 16546 21534 16558 21586
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 25666 21534 25678 21586
rect 25730 21534 25742 21586
rect 16158 21522 16210 21534
rect 10658 21422 10670 21474
rect 10722 21422 10734 21474
rect 21858 21422 21870 21474
rect 21922 21422 21934 21474
rect 25218 21422 25230 21474
rect 25282 21422 25294 21474
rect 15038 21362 15090 21374
rect 15038 21298 15090 21310
rect 16494 21362 16546 21374
rect 16494 21298 16546 21310
rect 16830 21362 16882 21374
rect 16830 21298 16882 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 14478 21026 14530 21038
rect 22990 21026 23042 21038
rect 20402 20974 20414 21026
rect 20466 20974 20478 21026
rect 21522 20974 21534 21026
rect 21586 20974 21598 21026
rect 14478 20962 14530 20974
rect 22990 20962 23042 20974
rect 24446 21026 24498 21038
rect 24446 20962 24498 20974
rect 15038 20914 15090 20926
rect 25454 20914 25506 20926
rect 40014 20914 40066 20926
rect 17154 20862 17166 20914
rect 17218 20862 17230 20914
rect 20066 20862 20078 20914
rect 20130 20862 20142 20914
rect 24210 20862 24222 20914
rect 24274 20862 24286 20914
rect 28578 20862 28590 20914
rect 28642 20862 28654 20914
rect 15038 20850 15090 20862
rect 25454 20850 25506 20862
rect 40014 20850 40066 20862
rect 15934 20802 15986 20814
rect 18062 20802 18114 20814
rect 14802 20750 14814 20802
rect 14866 20750 14878 20802
rect 17042 20750 17054 20802
rect 17106 20750 17118 20802
rect 15934 20738 15986 20750
rect 18062 20738 18114 20750
rect 18398 20802 18450 20814
rect 18398 20738 18450 20750
rect 18958 20802 19010 20814
rect 20302 20802 20354 20814
rect 19842 20750 19854 20802
rect 19906 20750 19918 20802
rect 18958 20738 19010 20750
rect 20302 20738 20354 20750
rect 21310 20802 21362 20814
rect 22878 20802 22930 20814
rect 29150 20802 29202 20814
rect 22306 20750 22318 20802
rect 22370 20750 22382 20802
rect 23538 20750 23550 20802
rect 23602 20750 23614 20802
rect 24098 20750 24110 20802
rect 24162 20750 24174 20802
rect 25666 20750 25678 20802
rect 25730 20750 25742 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 21310 20738 21362 20750
rect 22878 20738 22930 20750
rect 29150 20738 29202 20750
rect 17390 20690 17442 20702
rect 26450 20638 26462 20690
rect 26514 20638 26526 20690
rect 17390 20626 17442 20638
rect 14926 20578 14978 20590
rect 14926 20514 14978 20526
rect 15150 20578 15202 20590
rect 15150 20514 15202 20526
rect 15710 20578 15762 20590
rect 15710 20514 15762 20526
rect 15822 20578 15874 20590
rect 17714 20526 17726 20578
rect 17778 20526 17790 20578
rect 23762 20526 23774 20578
rect 23826 20526 23838 20578
rect 29474 20526 29486 20578
rect 29538 20526 29550 20578
rect 15822 20514 15874 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 24110 20242 24162 20254
rect 15474 20190 15486 20242
rect 15538 20190 15550 20242
rect 24110 20178 24162 20190
rect 26126 20242 26178 20254
rect 26126 20178 26178 20190
rect 11902 20130 11954 20142
rect 11902 20066 11954 20078
rect 14254 20130 14306 20142
rect 14254 20066 14306 20078
rect 17502 20130 17554 20142
rect 17502 20066 17554 20078
rect 17726 20130 17778 20142
rect 21422 20130 21474 20142
rect 18162 20078 18174 20130
rect 18226 20078 18238 20130
rect 17726 20066 17778 20078
rect 21422 20066 21474 20078
rect 22766 20130 22818 20142
rect 25790 20130 25842 20142
rect 24434 20078 24446 20130
rect 24498 20078 24510 20130
rect 22766 20066 22818 20078
rect 25790 20066 25842 20078
rect 14926 20018 14978 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 11666 19966 11678 20018
rect 11730 19966 11742 20018
rect 13906 19966 13918 20018
rect 13970 19966 13982 20018
rect 14926 19954 14978 19966
rect 15150 20018 15202 20030
rect 15934 20018 15986 20030
rect 20302 20018 20354 20030
rect 15586 19966 15598 20018
rect 15650 19966 15662 20018
rect 19954 19966 19966 20018
rect 20018 19966 20030 20018
rect 15150 19954 15202 19966
rect 15934 19954 15986 19966
rect 20302 19954 20354 19966
rect 22990 20018 23042 20030
rect 22990 19954 23042 19966
rect 26014 20018 26066 20030
rect 26014 19954 26066 19966
rect 26238 20018 26290 20030
rect 26238 19954 26290 19966
rect 26462 20018 26514 20030
rect 26462 19954 26514 19966
rect 26798 20018 26850 20030
rect 26798 19954 26850 19966
rect 27022 20018 27074 20030
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 27022 19954 27074 19966
rect 14142 19906 14194 19918
rect 26686 19906 26738 19918
rect 17378 19854 17390 19906
rect 17442 19854 17454 19906
rect 18610 19854 18622 19906
rect 18674 19854 18686 19906
rect 14142 19842 14194 19854
rect 26686 19842 26738 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 15374 19794 15426 19806
rect 15374 19730 15426 19742
rect 23214 19794 23266 19806
rect 23214 19730 23266 19742
rect 23438 19794 23490 19806
rect 23438 19730 23490 19742
rect 23886 19794 23938 19806
rect 23886 19730 23938 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 15038 19458 15090 19470
rect 15038 19394 15090 19406
rect 15486 19458 15538 19470
rect 23550 19458 23602 19470
rect 22306 19406 22318 19458
rect 22370 19406 22382 19458
rect 15486 19394 15538 19406
rect 23550 19394 23602 19406
rect 24894 19458 24946 19470
rect 24894 19394 24946 19406
rect 1934 19346 1986 19358
rect 25118 19346 25170 19358
rect 9986 19294 9998 19346
rect 10050 19294 10062 19346
rect 12114 19294 12126 19346
rect 12178 19294 12190 19346
rect 17602 19294 17614 19346
rect 17666 19294 17678 19346
rect 19618 19294 19630 19346
rect 19682 19294 19694 19346
rect 1934 19282 1986 19294
rect 25118 19282 25170 19294
rect 40014 19346 40066 19358
rect 40014 19282 40066 19294
rect 13582 19234 13634 19246
rect 14590 19234 14642 19246
rect 4274 19182 4286 19234
rect 4338 19182 4350 19234
rect 12898 19182 12910 19234
rect 12962 19182 12974 19234
rect 14354 19182 14366 19234
rect 14418 19182 14430 19234
rect 13582 19170 13634 19182
rect 14590 19170 14642 19182
rect 14814 19234 14866 19246
rect 22990 19234 23042 19246
rect 17266 19182 17278 19234
rect 17330 19182 17342 19234
rect 17826 19182 17838 19234
rect 17890 19182 17902 19234
rect 19394 19182 19406 19234
rect 19458 19182 19470 19234
rect 20514 19182 20526 19234
rect 20578 19182 20590 19234
rect 21970 19182 21982 19234
rect 22034 19182 22046 19234
rect 22530 19182 22542 19234
rect 22594 19182 22606 19234
rect 14814 19170 14866 19182
rect 22990 19170 23042 19182
rect 23102 19234 23154 19246
rect 23102 19170 23154 19182
rect 23326 19234 23378 19246
rect 23326 19170 23378 19182
rect 25454 19234 25506 19246
rect 25454 19170 25506 19182
rect 25566 19234 25618 19246
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 25566 19170 25618 19182
rect 15710 19122 15762 19134
rect 21758 19122 21810 19134
rect 16818 19070 16830 19122
rect 16882 19070 16894 19122
rect 19730 19070 19742 19122
rect 19794 19070 19806 19122
rect 20290 19070 20302 19122
rect 20354 19070 20366 19122
rect 15710 19058 15762 19070
rect 21758 19058 21810 19070
rect 14478 19010 14530 19022
rect 14478 18946 14530 18958
rect 15598 19010 15650 19022
rect 15598 18946 15650 18958
rect 22542 19010 22594 19022
rect 22542 18946 22594 18958
rect 23438 19010 23490 19022
rect 23438 18946 23490 18958
rect 25342 19010 25394 19022
rect 25342 18946 25394 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 19630 18674 19682 18686
rect 20626 18622 20638 18674
rect 20690 18622 20702 18674
rect 19630 18610 19682 18622
rect 17726 18562 17778 18574
rect 25790 18562 25842 18574
rect 16594 18510 16606 18562
rect 16658 18510 16670 18562
rect 18946 18510 18958 18562
rect 19010 18510 19022 18562
rect 19954 18510 19966 18562
rect 20018 18510 20030 18562
rect 22530 18510 22542 18562
rect 22594 18510 22606 18562
rect 17726 18498 17778 18510
rect 25790 18498 25842 18510
rect 26126 18562 26178 18574
rect 26126 18498 26178 18510
rect 26238 18562 26290 18574
rect 26238 18498 26290 18510
rect 15374 18450 15426 18462
rect 17838 18450 17890 18462
rect 14130 18398 14142 18450
rect 14194 18398 14206 18450
rect 14914 18398 14926 18450
rect 14978 18398 14990 18450
rect 16370 18398 16382 18450
rect 16434 18398 16446 18450
rect 15374 18386 15426 18398
rect 17838 18386 17890 18398
rect 18062 18450 18114 18462
rect 18622 18450 18674 18462
rect 18274 18398 18286 18450
rect 18338 18398 18350 18450
rect 18062 18386 18114 18398
rect 18622 18386 18674 18398
rect 20302 18450 20354 18462
rect 25230 18450 25282 18462
rect 21858 18398 21870 18450
rect 21922 18398 21934 18450
rect 20302 18386 20354 18398
rect 25230 18386 25282 18398
rect 25566 18450 25618 18462
rect 37874 18398 37886 18450
rect 37938 18398 37950 18450
rect 25566 18386 25618 18398
rect 25678 18338 25730 18350
rect 12002 18286 12014 18338
rect 12066 18286 12078 18338
rect 24658 18286 24670 18338
rect 24722 18286 24734 18338
rect 25678 18274 25730 18286
rect 26798 18338 26850 18350
rect 26798 18274 26850 18286
rect 26238 18226 26290 18238
rect 26238 18162 26290 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 16046 17890 16098 17902
rect 16046 17826 16098 17838
rect 1934 17778 1986 17790
rect 1934 17714 1986 17726
rect 16270 17778 16322 17790
rect 25006 17778 25058 17790
rect 40014 17778 40066 17790
rect 19058 17726 19070 17778
rect 19122 17726 19134 17778
rect 26114 17726 26126 17778
rect 26178 17726 26190 17778
rect 28242 17726 28254 17778
rect 28306 17726 28318 17778
rect 16270 17714 16322 17726
rect 25006 17714 25058 17726
rect 40014 17714 40066 17726
rect 22766 17666 22818 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 25330 17614 25342 17666
rect 25394 17614 25406 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 22766 17602 22818 17614
rect 19182 17554 19234 17566
rect 19182 17490 19234 17502
rect 19406 17554 19458 17566
rect 19406 17490 19458 17502
rect 19742 17554 19794 17566
rect 19742 17490 19794 17502
rect 20078 17554 20130 17566
rect 20078 17490 20130 17502
rect 20302 17554 20354 17566
rect 22418 17502 22430 17554
rect 22482 17502 22494 17554
rect 20302 17490 20354 17502
rect 19966 17442 20018 17454
rect 15698 17390 15710 17442
rect 15762 17390 15774 17442
rect 19966 17378 20018 17390
rect 20190 17442 20242 17454
rect 20190 17378 20242 17390
rect 24446 17442 24498 17454
rect 24446 17378 24498 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 15374 17106 15426 17118
rect 15374 17042 15426 17054
rect 16158 17106 16210 17118
rect 16158 17042 16210 17054
rect 16382 17106 16434 17118
rect 16382 17042 16434 17054
rect 16494 17106 16546 17118
rect 16494 17042 16546 17054
rect 21858 16942 21870 16994
rect 21922 16942 21934 16994
rect 27906 16942 27918 16994
rect 27970 16942 27982 16994
rect 15922 16830 15934 16882
rect 15986 16830 15998 16882
rect 19506 16830 19518 16882
rect 19570 16830 19582 16882
rect 27682 16830 27694 16882
rect 27746 16830 27758 16882
rect 15486 16770 15538 16782
rect 15486 16706 15538 16718
rect 16270 16770 16322 16782
rect 16270 16706 16322 16718
rect 15598 16658 15650 16670
rect 15598 16594 15650 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 24446 16322 24498 16334
rect 24446 16258 24498 16270
rect 16830 16210 16882 16222
rect 13458 16158 13470 16210
rect 13522 16158 13534 16210
rect 15586 16158 15598 16210
rect 15650 16158 15662 16210
rect 18610 16158 18622 16210
rect 18674 16158 18686 16210
rect 20738 16158 20750 16210
rect 20802 16158 20814 16210
rect 16830 16146 16882 16158
rect 16258 16046 16270 16098
rect 16322 16046 16334 16098
rect 17826 16046 17838 16098
rect 17890 16046 17902 16098
rect 21858 16046 21870 16098
rect 21922 16046 21934 16098
rect 21534 15986 21586 15998
rect 21534 15922 21586 15934
rect 21646 15874 21698 15886
rect 21646 15810 21698 15822
rect 22318 15874 22370 15886
rect 22318 15810 22370 15822
rect 24222 15874 24274 15886
rect 24222 15810 24274 15822
rect 24334 15874 24386 15886
rect 24334 15810 24386 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 20302 15538 20354 15550
rect 20302 15474 20354 15486
rect 20638 15538 20690 15550
rect 20638 15474 20690 15486
rect 23438 15538 23490 15550
rect 23438 15474 23490 15486
rect 25342 15538 25394 15550
rect 25342 15474 25394 15486
rect 25790 15538 25842 15550
rect 25790 15474 25842 15486
rect 17950 15426 18002 15438
rect 17950 15362 18002 15374
rect 19518 15426 19570 15438
rect 19518 15362 19570 15374
rect 20078 15426 20130 15438
rect 23214 15426 23266 15438
rect 21522 15374 21534 15426
rect 21586 15374 21598 15426
rect 20078 15362 20130 15374
rect 23214 15362 23266 15374
rect 16158 15314 16210 15326
rect 15586 15262 15598 15314
rect 15650 15262 15662 15314
rect 16158 15250 16210 15262
rect 16606 15314 16658 15326
rect 16606 15250 16658 15262
rect 16718 15314 16770 15326
rect 16718 15250 16770 15262
rect 17390 15314 17442 15326
rect 17390 15250 17442 15262
rect 17726 15314 17778 15326
rect 17726 15250 17778 15262
rect 20526 15314 20578 15326
rect 20526 15250 20578 15262
rect 21198 15314 21250 15326
rect 21198 15250 21250 15262
rect 23998 15314 24050 15326
rect 23998 15250 24050 15262
rect 24222 15314 24274 15326
rect 24222 15250 24274 15262
rect 15934 15202 15986 15214
rect 15934 15138 15986 15150
rect 16382 15202 16434 15214
rect 16382 15138 16434 15150
rect 17502 15202 17554 15214
rect 17502 15138 17554 15150
rect 19630 15202 19682 15214
rect 19630 15138 19682 15150
rect 19742 15202 19794 15214
rect 19742 15138 19794 15150
rect 20414 15202 20466 15214
rect 23538 15150 23550 15202
rect 23602 15150 23614 15202
rect 20414 15138 20466 15150
rect 15598 15090 15650 15102
rect 15598 15026 15650 15038
rect 23886 15090 23938 15102
rect 23886 15026 23938 15038
rect 24334 15090 24386 15102
rect 24334 15026 24386 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 18062 14754 18114 14766
rect 18062 14690 18114 14702
rect 18846 14642 18898 14654
rect 15586 14590 15598 14642
rect 15650 14590 15662 14642
rect 17714 14590 17726 14642
rect 17778 14590 17790 14642
rect 25106 14590 25118 14642
rect 25170 14590 25182 14642
rect 26226 14590 26238 14642
rect 26290 14590 26302 14642
rect 28354 14590 28366 14642
rect 28418 14590 28430 14642
rect 18846 14578 18898 14590
rect 14914 14478 14926 14530
rect 14978 14478 14990 14530
rect 18386 14478 18398 14530
rect 18450 14478 18462 14530
rect 22306 14478 22318 14530
rect 22370 14478 22382 14530
rect 25442 14478 25454 14530
rect 25506 14478 25518 14530
rect 22978 14366 22990 14418
rect 23042 14366 23054 14418
rect 18174 14306 18226 14318
rect 18174 14242 18226 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 17502 13970 17554 13982
rect 17502 13906 17554 13918
rect 23214 13970 23266 13982
rect 23214 13906 23266 13918
rect 25342 13970 25394 13982
rect 25342 13906 25394 13918
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 19954 13806 19966 13858
rect 20018 13806 20030 13858
rect 22878 13746 22930 13758
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 19282 13694 19294 13746
rect 19346 13694 19358 13746
rect 22878 13682 22930 13694
rect 23102 13746 23154 13758
rect 23314 13694 23326 13746
rect 23378 13694 23390 13746
rect 25554 13694 25566 13746
rect 25618 13694 25630 13746
rect 23102 13682 23154 13694
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 22082 13582 22094 13634
rect 22146 13582 22158 13634
rect 25230 13522 25282 13534
rect 25230 13458 25282 13470
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 22430 13074 22482 13086
rect 22430 13010 22482 13022
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 22318 5234 22370 5246
rect 22318 5170 22370 5182
rect 21298 5070 21310 5122
rect 21362 5070 21374 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 17378 4286 17390 4338
rect 17442 4286 17454 4338
rect 21074 4286 21086 4338
rect 21138 4286 21150 4338
rect 27906 4286 27918 4338
rect 27970 4286 27982 4338
rect 18398 4114 18450 4126
rect 18398 4050 18450 4062
rect 22094 4114 22146 4126
rect 22094 4050 22146 4062
rect 26014 4114 26066 4126
rect 26014 4050 26066 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 22430 3666 22482 3678
rect 22430 3602 22482 3614
rect 26126 3666 26178 3678
rect 26126 3602 26178 3614
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 21410 3502 21422 3554
rect 21474 3502 21486 3554
rect 25330 3502 25342 3554
rect 25394 3502 25406 3554
rect 17278 3330 17330 3342
rect 17278 3266 17330 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
rect 17266 1710 17278 1762
rect 17330 1759 17342 1762
rect 18162 1759 18174 1762
rect 17330 1713 18174 1759
rect 17330 1710 17342 1713
rect 18162 1710 18174 1713
rect 18226 1710 18238 1762
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18622 38222 18674 38274
rect 25566 38222 25618 38274
rect 17614 37998 17666 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 26798 37438 26850 37490
rect 25790 37214 25842 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 21422 28478 21474 28530
rect 17838 28366 17890 28418
rect 21310 28366 21362 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 15262 28030 15314 28082
rect 25342 28030 25394 28082
rect 14702 27918 14754 27970
rect 17950 27918 18002 27970
rect 18734 27918 18786 27970
rect 20862 27918 20914 27970
rect 23998 27918 24050 27970
rect 4286 27806 4338 27858
rect 14254 27806 14306 27858
rect 14478 27806 14530 27858
rect 14814 27806 14866 27858
rect 17390 27806 17442 27858
rect 17614 27806 17666 27858
rect 17838 27806 17890 27858
rect 18398 27806 18450 27858
rect 20190 27806 20242 27858
rect 23774 27806 23826 27858
rect 24110 27806 24162 27858
rect 25118 27806 25170 27858
rect 25454 27806 25506 27858
rect 11342 27694 11394 27746
rect 13470 27694 13522 27746
rect 16830 27694 16882 27746
rect 17726 27694 17778 27746
rect 22990 27694 23042 27746
rect 23438 27694 23490 27746
rect 1934 27582 1986 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 27470 27246 27522 27298
rect 1934 27134 1986 27186
rect 15374 27134 15426 27186
rect 17502 27134 17554 27186
rect 18622 27134 18674 27186
rect 20750 27134 20802 27186
rect 21646 27134 21698 27186
rect 23774 27134 23826 27186
rect 25902 27134 25954 27186
rect 40014 27134 40066 27186
rect 4286 27022 4338 27074
rect 14366 27022 14418 27074
rect 14590 27022 14642 27074
rect 17950 27022 18002 27074
rect 21310 27022 21362 27074
rect 21534 27022 21586 27074
rect 21758 27022 21810 27074
rect 21982 27022 22034 27074
rect 22990 27022 23042 27074
rect 27134 27022 27186 27074
rect 27582 27022 27634 27074
rect 37662 27022 37714 27074
rect 13918 26910 13970 26962
rect 26798 26910 26850 26962
rect 26910 26910 26962 26962
rect 13694 26798 13746 26850
rect 13806 26798 13858 26850
rect 26350 26798 26402 26850
rect 27470 26798 27522 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 15150 26462 15202 26514
rect 15822 26462 15874 26514
rect 20974 26462 21026 26514
rect 21982 26462 22034 26514
rect 24670 26462 24722 26514
rect 13918 26350 13970 26402
rect 16046 26350 16098 26402
rect 16494 26350 16546 26402
rect 18510 26350 18562 26402
rect 18846 26350 18898 26402
rect 18958 26350 19010 26402
rect 23662 26350 23714 26402
rect 26238 26350 26290 26402
rect 14590 26238 14642 26290
rect 14926 26238 14978 26290
rect 15262 26238 15314 26290
rect 16158 26238 16210 26290
rect 16830 26238 16882 26290
rect 17838 26238 17890 26290
rect 19182 26238 19234 26290
rect 19518 26238 19570 26290
rect 21758 26238 21810 26290
rect 23550 26238 23602 26290
rect 23886 26238 23938 26290
rect 25454 26238 25506 26290
rect 11790 26126 11842 26178
rect 17614 26126 17666 26178
rect 28366 26126 28418 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 17614 25678 17666 25730
rect 13582 25566 13634 25618
rect 14926 25566 14978 25618
rect 19294 25566 19346 25618
rect 22878 25566 22930 25618
rect 25006 25566 25058 25618
rect 26238 25566 26290 25618
rect 40014 25566 40066 25618
rect 13470 25454 13522 25506
rect 14142 25454 14194 25506
rect 16158 25454 16210 25506
rect 18174 25454 18226 25506
rect 19966 25454 20018 25506
rect 25678 25454 25730 25506
rect 27022 25454 27074 25506
rect 37662 25454 37714 25506
rect 16382 25342 16434 25394
rect 16494 25342 16546 25394
rect 17726 25342 17778 25394
rect 17950 25342 18002 25394
rect 19182 25342 19234 25394
rect 19406 25342 19458 25394
rect 27134 25342 27186 25394
rect 13694 25230 13746 25282
rect 16942 25230 16994 25282
rect 17390 25230 17442 25282
rect 19742 25230 19794 25282
rect 27358 25230 27410 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 18286 24894 18338 24946
rect 18622 24894 18674 24946
rect 25454 24894 25506 24946
rect 22990 24782 23042 24834
rect 19518 24670 19570 24722
rect 25790 24670 25842 24722
rect 26574 24558 26626 24610
rect 28702 24558 28754 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 23662 24110 23714 24162
rect 26462 24110 26514 24162
rect 1934 23998 1986 24050
rect 16382 23998 16434 24050
rect 17614 23998 17666 24050
rect 21870 23998 21922 24050
rect 24782 23998 24834 24050
rect 25342 23998 25394 24050
rect 4286 23886 4338 23938
rect 13582 23886 13634 23938
rect 16830 23886 16882 23938
rect 20638 23886 20690 23938
rect 21422 23886 21474 23938
rect 22318 23886 22370 23938
rect 24334 23886 24386 23938
rect 26574 23886 26626 23938
rect 14254 23774 14306 23826
rect 20302 23774 20354 23826
rect 22878 23774 22930 23826
rect 23214 23774 23266 23826
rect 23774 23774 23826 23826
rect 17166 23662 17218 23714
rect 20638 23662 20690 23714
rect 21310 23662 21362 23714
rect 23662 23662 23714 23714
rect 26462 23662 26514 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 14366 23326 14418 23378
rect 17726 23326 17778 23378
rect 18958 23326 19010 23378
rect 21870 23326 21922 23378
rect 24222 23326 24274 23378
rect 18622 23214 18674 23266
rect 22990 23214 23042 23266
rect 13694 23102 13746 23154
rect 14478 23102 14530 23154
rect 15374 23102 15426 23154
rect 20862 23102 20914 23154
rect 21758 23102 21810 23154
rect 22766 23102 22818 23154
rect 23662 23102 23714 23154
rect 24446 23102 24498 23154
rect 28254 23102 28306 23154
rect 10894 22990 10946 23042
rect 13022 22990 13074 23042
rect 15710 22990 15762 23042
rect 18286 22990 18338 23042
rect 19630 22990 19682 23042
rect 19966 22990 20018 23042
rect 20414 22990 20466 23042
rect 21534 22990 21586 23042
rect 25454 22990 25506 23042
rect 27582 22990 27634 23042
rect 14366 22878 14418 22930
rect 15150 22878 15202 22930
rect 15262 22878 15314 22930
rect 15934 22878 15986 22930
rect 22430 22878 22482 22930
rect 23326 22878 23378 22930
rect 23438 22878 23490 22930
rect 23774 22878 23826 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 17278 22542 17330 22594
rect 17950 22542 18002 22594
rect 25230 22542 25282 22594
rect 26350 22542 26402 22594
rect 1934 22430 1986 22482
rect 14030 22430 14082 22482
rect 19294 22430 19346 22482
rect 4286 22318 4338 22370
rect 17166 22318 17218 22370
rect 17726 22318 17778 22370
rect 18286 22318 18338 22370
rect 20190 22318 20242 22370
rect 20750 22318 20802 22370
rect 22878 22318 22930 22370
rect 24782 22318 24834 22370
rect 25118 22318 25170 22370
rect 25678 22318 25730 22370
rect 18510 22206 18562 22258
rect 22094 22206 22146 22258
rect 23102 22206 23154 22258
rect 24894 22206 24946 22258
rect 26238 22206 26290 22258
rect 17614 22094 17666 22146
rect 18846 22094 18898 22146
rect 19854 22094 19906 22146
rect 25230 22094 25282 22146
rect 25790 22094 25842 22146
rect 26014 22094 26066 22146
rect 26350 22094 26402 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14030 21758 14082 21810
rect 14702 21758 14754 21810
rect 12798 21646 12850 21698
rect 15262 21646 15314 21698
rect 15822 21646 15874 21698
rect 18174 21646 18226 21698
rect 18510 21646 18562 21698
rect 19070 21646 19122 21698
rect 25566 21646 25618 21698
rect 40238 21646 40290 21698
rect 13582 21534 13634 21586
rect 14926 21534 14978 21586
rect 15486 21534 15538 21586
rect 16158 21534 16210 21586
rect 16494 21534 16546 21586
rect 17838 21534 17890 21586
rect 19406 21534 19458 21586
rect 25678 21534 25730 21586
rect 10670 21422 10722 21474
rect 21870 21422 21922 21474
rect 25230 21422 25282 21474
rect 15038 21310 15090 21362
rect 16494 21310 16546 21362
rect 16830 21310 16882 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 14478 20974 14530 21026
rect 20414 20974 20466 21026
rect 21534 20974 21586 21026
rect 22990 20974 23042 21026
rect 24446 20974 24498 21026
rect 15038 20862 15090 20914
rect 17166 20862 17218 20914
rect 20078 20862 20130 20914
rect 24222 20862 24274 20914
rect 25454 20862 25506 20914
rect 28590 20862 28642 20914
rect 40014 20862 40066 20914
rect 14814 20750 14866 20802
rect 15934 20750 15986 20802
rect 17054 20750 17106 20802
rect 18062 20750 18114 20802
rect 18398 20750 18450 20802
rect 18958 20750 19010 20802
rect 19854 20750 19906 20802
rect 20302 20750 20354 20802
rect 21310 20750 21362 20802
rect 22318 20750 22370 20802
rect 22878 20750 22930 20802
rect 23550 20750 23602 20802
rect 24110 20750 24162 20802
rect 25678 20750 25730 20802
rect 29150 20750 29202 20802
rect 37662 20750 37714 20802
rect 17390 20638 17442 20690
rect 26462 20638 26514 20690
rect 14926 20526 14978 20578
rect 15150 20526 15202 20578
rect 15710 20526 15762 20578
rect 15822 20526 15874 20578
rect 17726 20526 17778 20578
rect 23774 20526 23826 20578
rect 29486 20526 29538 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 15486 20190 15538 20242
rect 24110 20190 24162 20242
rect 26126 20190 26178 20242
rect 11902 20078 11954 20130
rect 14254 20078 14306 20130
rect 17502 20078 17554 20130
rect 17726 20078 17778 20130
rect 18174 20078 18226 20130
rect 21422 20078 21474 20130
rect 22766 20078 22818 20130
rect 24446 20078 24498 20130
rect 25790 20078 25842 20130
rect 4286 19966 4338 20018
rect 11678 19966 11730 20018
rect 13918 19966 13970 20018
rect 14926 19966 14978 20018
rect 15150 19966 15202 20018
rect 15598 19966 15650 20018
rect 15934 19966 15986 20018
rect 19966 19966 20018 20018
rect 20302 19966 20354 20018
rect 22990 19966 23042 20018
rect 26014 19966 26066 20018
rect 26238 19966 26290 20018
rect 26462 19966 26514 20018
rect 26798 19966 26850 20018
rect 27022 19966 27074 20018
rect 37662 19966 37714 20018
rect 14142 19854 14194 19906
rect 17390 19854 17442 19906
rect 18622 19854 18674 19906
rect 26686 19854 26738 19906
rect 1934 19742 1986 19794
rect 15374 19742 15426 19794
rect 23214 19742 23266 19794
rect 23438 19742 23490 19794
rect 23886 19742 23938 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15038 19406 15090 19458
rect 15486 19406 15538 19458
rect 22318 19406 22370 19458
rect 23550 19406 23602 19458
rect 24894 19406 24946 19458
rect 1934 19294 1986 19346
rect 9998 19294 10050 19346
rect 12126 19294 12178 19346
rect 17614 19294 17666 19346
rect 19630 19294 19682 19346
rect 25118 19294 25170 19346
rect 40014 19294 40066 19346
rect 4286 19182 4338 19234
rect 12910 19182 12962 19234
rect 13582 19182 13634 19234
rect 14366 19182 14418 19234
rect 14590 19182 14642 19234
rect 14814 19182 14866 19234
rect 17278 19182 17330 19234
rect 17838 19182 17890 19234
rect 19406 19182 19458 19234
rect 20526 19182 20578 19234
rect 21982 19182 22034 19234
rect 22542 19182 22594 19234
rect 22990 19182 23042 19234
rect 23102 19182 23154 19234
rect 23326 19182 23378 19234
rect 25454 19182 25506 19234
rect 25566 19182 25618 19234
rect 37662 19182 37714 19234
rect 15710 19070 15762 19122
rect 16830 19070 16882 19122
rect 19742 19070 19794 19122
rect 20302 19070 20354 19122
rect 21758 19070 21810 19122
rect 14478 18958 14530 19010
rect 15598 18958 15650 19010
rect 22542 18958 22594 19010
rect 23438 18958 23490 19010
rect 25342 18958 25394 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 19630 18622 19682 18674
rect 20638 18622 20690 18674
rect 16606 18510 16658 18562
rect 17726 18510 17778 18562
rect 18958 18510 19010 18562
rect 19966 18510 20018 18562
rect 22542 18510 22594 18562
rect 25790 18510 25842 18562
rect 26126 18510 26178 18562
rect 26238 18510 26290 18562
rect 14142 18398 14194 18450
rect 14926 18398 14978 18450
rect 15374 18398 15426 18450
rect 16382 18398 16434 18450
rect 17838 18398 17890 18450
rect 18062 18398 18114 18450
rect 18286 18398 18338 18450
rect 18622 18398 18674 18450
rect 20302 18398 20354 18450
rect 21870 18398 21922 18450
rect 25230 18398 25282 18450
rect 25566 18398 25618 18450
rect 37886 18398 37938 18450
rect 12014 18286 12066 18338
rect 24670 18286 24722 18338
rect 25678 18286 25730 18338
rect 26798 18286 26850 18338
rect 26238 18174 26290 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 16046 17838 16098 17890
rect 1934 17726 1986 17778
rect 16270 17726 16322 17778
rect 19070 17726 19122 17778
rect 25006 17726 25058 17778
rect 26126 17726 26178 17778
rect 28254 17726 28306 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 22766 17614 22818 17666
rect 25342 17614 25394 17666
rect 37662 17614 37714 17666
rect 19182 17502 19234 17554
rect 19406 17502 19458 17554
rect 19742 17502 19794 17554
rect 20078 17502 20130 17554
rect 20302 17502 20354 17554
rect 22430 17502 22482 17554
rect 15710 17390 15762 17442
rect 19966 17390 20018 17442
rect 20190 17390 20242 17442
rect 24446 17390 24498 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 15374 17054 15426 17106
rect 16158 17054 16210 17106
rect 16382 17054 16434 17106
rect 16494 17054 16546 17106
rect 21870 16942 21922 16994
rect 27918 16942 27970 16994
rect 15934 16830 15986 16882
rect 19518 16830 19570 16882
rect 27694 16830 27746 16882
rect 15486 16718 15538 16770
rect 16270 16718 16322 16770
rect 15598 16606 15650 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 24446 16270 24498 16322
rect 13470 16158 13522 16210
rect 15598 16158 15650 16210
rect 16830 16158 16882 16210
rect 18622 16158 18674 16210
rect 20750 16158 20802 16210
rect 16270 16046 16322 16098
rect 17838 16046 17890 16098
rect 21870 16046 21922 16098
rect 21534 15934 21586 15986
rect 21646 15822 21698 15874
rect 22318 15822 22370 15874
rect 24222 15822 24274 15874
rect 24334 15822 24386 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 20302 15486 20354 15538
rect 20638 15486 20690 15538
rect 23438 15486 23490 15538
rect 25342 15486 25394 15538
rect 25790 15486 25842 15538
rect 17950 15374 18002 15426
rect 19518 15374 19570 15426
rect 20078 15374 20130 15426
rect 21534 15374 21586 15426
rect 23214 15374 23266 15426
rect 15598 15262 15650 15314
rect 16158 15262 16210 15314
rect 16606 15262 16658 15314
rect 16718 15262 16770 15314
rect 17390 15262 17442 15314
rect 17726 15262 17778 15314
rect 20526 15262 20578 15314
rect 21198 15262 21250 15314
rect 23998 15262 24050 15314
rect 24222 15262 24274 15314
rect 15934 15150 15986 15202
rect 16382 15150 16434 15202
rect 17502 15150 17554 15202
rect 19630 15150 19682 15202
rect 19742 15150 19794 15202
rect 20414 15150 20466 15202
rect 23550 15150 23602 15202
rect 15598 15038 15650 15090
rect 23886 15038 23938 15090
rect 24334 15038 24386 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 18062 14702 18114 14754
rect 15598 14590 15650 14642
rect 17726 14590 17778 14642
rect 18846 14590 18898 14642
rect 25118 14590 25170 14642
rect 26238 14590 26290 14642
rect 28366 14590 28418 14642
rect 14926 14478 14978 14530
rect 18398 14478 18450 14530
rect 22318 14478 22370 14530
rect 25454 14478 25506 14530
rect 22990 14366 23042 14418
rect 18174 14254 18226 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17502 13918 17554 13970
rect 23214 13918 23266 13970
rect 25342 13918 25394 13970
rect 14702 13806 14754 13858
rect 19966 13806 20018 13858
rect 14030 13694 14082 13746
rect 19294 13694 19346 13746
rect 22878 13694 22930 13746
rect 23102 13694 23154 13746
rect 23326 13694 23378 13746
rect 25566 13694 25618 13746
rect 16830 13582 16882 13634
rect 22094 13582 22146 13634
rect 25230 13470 25282 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 22430 13022 22482 13074
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 22318 5182 22370 5234
rect 21310 5070 21362 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 17390 4286 17442 4338
rect 21086 4286 21138 4338
rect 27918 4286 27970 4338
rect 18398 4062 18450 4114
rect 22094 4062 22146 4114
rect 26014 4062 26066 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 22430 3614 22482 3666
rect 26126 3614 26178 3666
rect 17614 3502 17666 3554
rect 21422 3502 21474 3554
rect 25342 3502 25394 3554
rect 17278 3278 17330 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 17278 1710 17330 1762
rect 18174 1710 18226 1762
<< metal2 >>
rect 18144 41200 18256 42000
rect 22848 41200 22960 42000
rect 25536 41200 25648 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 18172 38276 18228 41200
rect 18620 38276 18676 38286
rect 18172 38274 18676 38276
rect 18172 38222 18622 38274
rect 18674 38222 18676 38274
rect 18172 38220 18676 38222
rect 18620 38210 18676 38220
rect 22876 38276 22932 41200
rect 25564 38612 25620 41200
rect 25564 38546 25620 38556
rect 26796 38612 26852 38622
rect 22876 38210 22932 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 17612 38050 17668 38062
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 17612 31948 17668 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 17500 31892 17668 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 14588 28084 14644 28094
rect 14252 28028 14588 28084
rect 4284 27860 4340 27870
rect 4284 27766 4340 27804
rect 11788 27860 11844 27870
rect 11340 27746 11396 27758
rect 11340 27694 11342 27746
rect 11394 27694 11396 27746
rect 1932 27636 1988 27646
rect 1932 27542 1988 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 27188 1988 27198
rect 1932 27094 1988 27132
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 11340 27076 11396 27694
rect 11340 27010 11396 27020
rect 4956 26292 5012 26302
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 4284 23938 4340 23950
rect 4284 23886 4286 23938
rect 4338 23886 4340 23938
rect 4284 23044 4340 23886
rect 4284 22978 4340 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 1932 22482 1988 22494
rect 1932 22430 1934 22482
rect 1986 22430 1988 22482
rect 1932 21588 1988 22430
rect 1932 21522 1988 21532
rect 4284 22370 4340 22382
rect 4284 22318 4286 22370
rect 4338 22318 4340 22370
rect 4284 21476 4340 22318
rect 4956 22148 5012 26236
rect 11788 26178 11844 27804
rect 14252 27858 14308 28028
rect 14252 27806 14254 27858
rect 14306 27806 14308 27858
rect 14252 27794 14308 27806
rect 14476 27858 14532 27870
rect 14476 27806 14478 27858
rect 14530 27806 14532 27858
rect 13468 27748 13524 27758
rect 13468 27746 13636 27748
rect 13468 27694 13470 27746
rect 13522 27694 13636 27746
rect 13468 27692 13636 27694
rect 13468 27682 13524 27692
rect 11788 26126 11790 26178
rect 11842 26126 11844 26178
rect 11788 26114 11844 26126
rect 13580 25618 13636 27692
rect 14364 27076 14420 27086
rect 14476 27076 14532 27806
rect 14364 27074 14532 27076
rect 14364 27022 14366 27074
rect 14418 27022 14532 27074
rect 14364 27020 14532 27022
rect 14588 27076 14644 28028
rect 15260 28084 15316 28094
rect 15260 27990 15316 28028
rect 14700 27970 14756 27982
rect 14700 27918 14702 27970
rect 14754 27918 14756 27970
rect 14700 27860 14756 27918
rect 16940 27972 16996 27982
rect 14700 27794 14756 27804
rect 14812 27860 14868 27870
rect 15820 27860 15876 27870
rect 14812 27858 15092 27860
rect 14812 27806 14814 27858
rect 14866 27806 15092 27858
rect 14812 27804 15092 27806
rect 14812 27794 14868 27804
rect 14588 27074 14756 27076
rect 14588 27022 14590 27074
rect 14642 27022 14756 27074
rect 14588 27020 14756 27022
rect 14364 27010 14420 27020
rect 14588 27010 14644 27020
rect 13916 26964 13972 26974
rect 13916 26962 14084 26964
rect 13916 26910 13918 26962
rect 13970 26910 14084 26962
rect 13916 26908 14084 26910
rect 13916 26898 13972 26908
rect 13580 25566 13582 25618
rect 13634 25566 13636 25618
rect 13580 25554 13636 25566
rect 13692 26850 13748 26862
rect 13692 26798 13694 26850
rect 13746 26798 13748 26850
rect 13468 25508 13524 25518
rect 13468 25414 13524 25452
rect 13692 25508 13748 26798
rect 13804 26850 13860 26862
rect 13804 26798 13806 26850
rect 13858 26798 13860 26850
rect 13804 26404 13860 26798
rect 13916 26404 13972 26414
rect 13804 26402 13972 26404
rect 13804 26350 13918 26402
rect 13970 26350 13972 26402
rect 13804 26348 13972 26350
rect 13916 26338 13972 26348
rect 14028 26404 14084 26908
rect 14700 26908 14756 27020
rect 14700 26852 14868 26908
rect 14028 26338 14084 26348
rect 14252 26292 14308 26302
rect 13692 25442 13748 25452
rect 14140 26236 14252 26292
rect 14140 25506 14196 26236
rect 14252 26226 14308 26236
rect 14588 26290 14644 26302
rect 14588 26238 14590 26290
rect 14642 26238 14644 26290
rect 14588 26180 14644 26238
rect 14812 26180 14868 26852
rect 14924 26292 14980 26302
rect 15036 26292 15092 27804
rect 15372 27188 15428 27198
rect 15372 27094 15428 27132
rect 15148 27076 15204 27086
rect 15148 26514 15204 27020
rect 15148 26462 15150 26514
rect 15202 26462 15204 26514
rect 15148 26450 15204 26462
rect 15820 26514 15876 27804
rect 16828 27748 16884 27758
rect 16940 27748 16996 27916
rect 17388 27860 17444 27870
rect 17388 27766 17444 27804
rect 16828 27746 16996 27748
rect 16828 27694 16830 27746
rect 16882 27694 16996 27746
rect 16828 27692 16996 27694
rect 16828 27682 16884 27692
rect 16044 27076 16100 27086
rect 15820 26462 15822 26514
rect 15874 26462 15876 26514
rect 15820 26450 15876 26462
rect 15932 27020 16044 27076
rect 15372 26404 15428 26414
rect 15260 26292 15316 26302
rect 15036 26290 15316 26292
rect 15036 26238 15262 26290
rect 15314 26238 15316 26290
rect 15036 26236 15316 26238
rect 14924 26198 14980 26236
rect 14588 26124 14868 26180
rect 14812 26068 14868 26124
rect 15260 26068 15316 26236
rect 14812 26012 14980 26068
rect 14140 25454 14142 25506
rect 14194 25454 14196 25506
rect 14140 25442 14196 25454
rect 14924 25618 14980 26012
rect 14924 25566 14926 25618
rect 14978 25566 14980 25618
rect 13692 25284 13748 25294
rect 13692 25282 13860 25284
rect 13692 25230 13694 25282
rect 13746 25230 13860 25282
rect 13692 25228 13860 25230
rect 13692 25218 13748 25228
rect 13580 24052 13636 24062
rect 13580 23940 13636 23996
rect 13580 23938 13748 23940
rect 13580 23886 13582 23938
rect 13634 23886 13748 23938
rect 13580 23884 13748 23886
rect 13580 23874 13636 23884
rect 10892 23380 10948 23390
rect 10892 23044 10948 23324
rect 13692 23156 13748 23884
rect 13804 23828 13860 25228
rect 14924 24052 14980 25566
rect 14924 23986 14980 23996
rect 14252 23828 14308 23838
rect 13804 23826 14308 23828
rect 13804 23774 14254 23826
rect 14306 23774 14308 23826
rect 13804 23772 14308 23774
rect 14252 23492 14308 23772
rect 14252 23426 14308 23436
rect 15036 23492 15092 23502
rect 14364 23380 14420 23390
rect 14364 23286 14420 23324
rect 14476 23156 14532 23166
rect 13692 23154 14084 23156
rect 13692 23102 13694 23154
rect 13746 23102 14084 23154
rect 13692 23100 14084 23102
rect 13692 23090 13748 23100
rect 10892 22950 10948 22988
rect 13020 23044 13076 23054
rect 13020 22950 13076 22988
rect 4956 22082 5012 22092
rect 14028 22482 14084 23100
rect 14476 23062 14532 23100
rect 14364 22932 14420 22942
rect 14364 22838 14420 22876
rect 14028 22430 14030 22482
rect 14082 22430 14084 22482
rect 12796 21812 12852 21822
rect 14028 21812 14084 22430
rect 14812 21924 14868 21934
rect 12796 21698 12852 21756
rect 12796 21646 12798 21698
rect 12850 21646 12852 21698
rect 12796 21634 12852 21646
rect 13580 21810 14084 21812
rect 13580 21758 14030 21810
rect 14082 21758 14084 21810
rect 13580 21756 14084 21758
rect 13580 21586 13636 21756
rect 14028 21746 14084 21756
rect 14700 21812 14756 21822
rect 14700 21718 14756 21756
rect 13580 21534 13582 21586
rect 13634 21534 13636 21586
rect 13580 21522 13636 21534
rect 4284 21410 4340 21420
rect 10668 21476 10724 21486
rect 10668 21382 10724 21420
rect 14476 21476 14532 21486
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 14476 21026 14532 21420
rect 14476 20974 14478 21026
rect 14530 20974 14532 21026
rect 14476 20962 14532 20974
rect 14812 20804 14868 21868
rect 15036 21812 15092 23436
rect 15260 23492 15316 26012
rect 15260 23426 15316 23436
rect 15372 23154 15428 26348
rect 15932 23156 15988 27020
rect 16044 27010 16100 27020
rect 16044 26404 16100 26414
rect 16044 26310 16100 26348
rect 16492 26404 16548 26414
rect 16492 26310 16548 26348
rect 16156 26292 16212 26302
rect 16828 26292 16884 26302
rect 16156 26290 16324 26292
rect 16156 26238 16158 26290
rect 16210 26238 16324 26290
rect 16156 26236 16324 26238
rect 16156 26226 16212 26236
rect 16156 25508 16212 25518
rect 16156 25414 16212 25452
rect 15372 23102 15374 23154
rect 15426 23102 15428 23154
rect 15260 23044 15316 23054
rect 15148 22932 15204 22942
rect 15148 22838 15204 22876
rect 15260 22930 15316 22988
rect 15260 22878 15262 22930
rect 15314 22878 15316 22930
rect 15260 22866 15316 22878
rect 15260 22036 15316 22046
rect 15036 21746 15092 21756
rect 15148 21980 15260 22036
rect 14924 21586 14980 21598
rect 14924 21534 14926 21586
rect 14978 21534 14980 21586
rect 14924 20916 14980 21534
rect 14924 20850 14980 20860
rect 15036 21362 15092 21374
rect 15036 21310 15038 21362
rect 15090 21310 15092 21362
rect 15036 20914 15092 21310
rect 15148 21364 15204 21980
rect 15260 21970 15316 21980
rect 15260 21812 15316 21822
rect 15260 21698 15316 21756
rect 15260 21646 15262 21698
rect 15314 21646 15316 21698
rect 15260 21634 15316 21646
rect 15148 21308 15316 21364
rect 15036 20862 15038 20914
rect 15090 20862 15092 20914
rect 15036 20850 15092 20862
rect 14252 20802 14868 20804
rect 14252 20750 14814 20802
rect 14866 20750 14868 20802
rect 14252 20748 14868 20750
rect 11900 20132 11956 20142
rect 11900 20130 12180 20132
rect 11900 20078 11902 20130
rect 11954 20078 12180 20130
rect 11900 20076 12180 20078
rect 11900 20066 11956 20076
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 9996 20020 10052 20030
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1932 19346 1988 19358
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 18900 1988 19294
rect 9996 19346 10052 19964
rect 11676 20018 11732 20030
rect 11676 19966 11678 20018
rect 11730 19966 11732 20018
rect 11676 19572 11732 19966
rect 11676 19506 11732 19516
rect 12012 19684 12068 19694
rect 9996 19294 9998 19346
rect 10050 19294 10052 19346
rect 9996 19282 10052 19294
rect 4284 19236 4340 19246
rect 4284 19142 4340 19180
rect 12012 19236 12068 19628
rect 12124 19346 12180 20076
rect 14252 20130 14308 20748
rect 14812 20738 14868 20748
rect 14924 20580 14980 20590
rect 14924 20486 14980 20524
rect 15148 20578 15204 20590
rect 15148 20526 15150 20578
rect 15202 20526 15204 20578
rect 15148 20244 15204 20526
rect 15148 20178 15204 20188
rect 14252 20078 14254 20130
rect 14306 20078 14308 20130
rect 14252 20066 14308 20078
rect 13916 20020 13972 20030
rect 13916 19926 13972 19964
rect 14924 20018 14980 20030
rect 14924 19966 14926 20018
rect 14978 19966 14980 20018
rect 12124 19294 12126 19346
rect 12178 19294 12180 19346
rect 12124 19282 12180 19294
rect 14140 19906 14196 19918
rect 14140 19854 14142 19906
rect 14194 19854 14196 19906
rect 1932 18834 1988 18844
rect 12012 18338 12068 19180
rect 12908 19236 12964 19246
rect 12908 19142 12964 19180
rect 13580 19236 13636 19246
rect 14140 19236 14196 19854
rect 14924 19684 14980 19966
rect 15148 20020 15204 20030
rect 15260 20020 15316 21308
rect 15372 20468 15428 23102
rect 15820 23100 15988 23156
rect 16268 25172 16324 26236
rect 16828 26198 16884 26236
rect 16380 26180 16436 26190
rect 16380 25394 16436 26124
rect 16380 25342 16382 25394
rect 16434 25342 16436 25394
rect 16380 25330 16436 25342
rect 16492 25394 16548 25406
rect 16492 25342 16494 25394
rect 16546 25342 16548 25394
rect 16492 25284 16548 25342
rect 16940 25284 16996 27692
rect 17500 27186 17556 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 21420 28532 21476 28542
rect 21420 28530 21700 28532
rect 21420 28478 21422 28530
rect 21474 28478 21700 28530
rect 21420 28476 21700 28478
rect 21420 28466 21476 28476
rect 17836 28418 17892 28430
rect 21308 28420 21364 28430
rect 17836 28366 17838 28418
rect 17890 28366 17892 28418
rect 17836 28196 17892 28366
rect 20860 28418 21364 28420
rect 20860 28366 21310 28418
rect 21362 28366 21364 28418
rect 20860 28364 21364 28366
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 17836 28140 18116 28196
rect 19836 28186 20100 28196
rect 17836 28084 17892 28140
rect 17836 28018 17892 28028
rect 17948 27972 18004 27982
rect 17948 27878 18004 27916
rect 17500 27134 17502 27186
rect 17554 27134 17556 27186
rect 17500 25396 17556 27134
rect 17612 27858 17668 27870
rect 17612 27806 17614 27858
rect 17666 27806 17668 27858
rect 17612 26908 17668 27806
rect 17836 27858 17892 27870
rect 17836 27806 17838 27858
rect 17890 27806 17892 27858
rect 17724 27746 17780 27758
rect 17724 27694 17726 27746
rect 17778 27694 17780 27746
rect 17724 27188 17780 27694
rect 17724 27122 17780 27132
rect 17612 26852 17780 26908
rect 17612 26180 17668 26190
rect 17612 26086 17668 26124
rect 17612 25732 17668 25742
rect 17724 25732 17780 26852
rect 17836 26516 17892 27806
rect 17948 27076 18004 27086
rect 18060 27076 18116 28140
rect 18732 27970 18788 27982
rect 18732 27918 18734 27970
rect 18786 27918 18788 27970
rect 17948 27074 18116 27076
rect 17948 27022 17950 27074
rect 18002 27022 18116 27074
rect 17948 27020 18116 27022
rect 18396 27858 18452 27870
rect 18396 27806 18398 27858
rect 18450 27806 18452 27858
rect 17948 26964 18004 27020
rect 17948 26898 18004 26908
rect 17836 26460 18004 26516
rect 17612 25730 17780 25732
rect 17612 25678 17614 25730
rect 17666 25678 17780 25730
rect 17612 25676 17780 25678
rect 17836 26292 17892 26302
rect 17612 25666 17668 25676
rect 17724 25396 17780 25406
rect 17500 25394 17780 25396
rect 17500 25342 17726 25394
rect 17778 25342 17780 25394
rect 17500 25340 17780 25342
rect 17724 25330 17780 25340
rect 17388 25284 17444 25294
rect 16492 25282 17444 25284
rect 16492 25230 16942 25282
rect 16994 25230 17390 25282
rect 17442 25230 17444 25282
rect 16492 25228 17444 25230
rect 16492 25172 16548 25228
rect 16940 25218 16996 25228
rect 17388 25218 17444 25228
rect 16268 25116 16548 25172
rect 15708 23044 15764 23054
rect 15708 22950 15764 22988
rect 15820 21698 15876 23100
rect 15932 22930 15988 22942
rect 15932 22878 15934 22930
rect 15986 22878 15988 22930
rect 15932 22820 15988 22878
rect 15932 22754 15988 22764
rect 15820 21646 15822 21698
rect 15874 21646 15876 21698
rect 15484 21586 15540 21598
rect 15484 21534 15486 21586
rect 15538 21534 15540 21586
rect 15484 21364 15540 21534
rect 15820 21588 15876 21646
rect 15820 21532 16100 21588
rect 15708 21364 15764 21374
rect 15484 21308 15708 21364
rect 15708 21298 15764 21308
rect 15932 20804 15988 20842
rect 15932 20738 15988 20748
rect 15708 20580 15764 20590
rect 15708 20486 15764 20524
rect 15820 20578 15876 20590
rect 15820 20526 15822 20578
rect 15874 20526 15876 20578
rect 15596 20468 15652 20478
rect 15372 20412 15596 20468
rect 15596 20402 15652 20412
rect 15148 20018 15316 20020
rect 15148 19966 15150 20018
rect 15202 19966 15316 20018
rect 15148 19964 15316 19966
rect 15484 20242 15540 20254
rect 15820 20244 15876 20526
rect 15484 20190 15486 20242
rect 15538 20190 15540 20242
rect 15148 19954 15204 19964
rect 14924 19618 14980 19628
rect 15372 19794 15428 19806
rect 15372 19742 15374 19794
rect 15426 19742 15428 19794
rect 14476 19572 14532 19582
rect 14364 19236 14420 19246
rect 14140 19234 14420 19236
rect 14140 19182 14366 19234
rect 14418 19182 14420 19234
rect 14140 19180 14420 19182
rect 13580 19142 13636 19180
rect 14364 19170 14420 19180
rect 14140 19012 14196 19022
rect 14140 18450 14196 18956
rect 14476 19010 14532 19516
rect 15036 19460 15092 19470
rect 15036 19366 15092 19404
rect 14588 19348 14644 19358
rect 14588 19234 14644 19292
rect 14588 19182 14590 19234
rect 14642 19182 14644 19234
rect 14588 19170 14644 19182
rect 14812 19234 14868 19246
rect 14812 19182 14814 19234
rect 14866 19182 14868 19234
rect 14476 18958 14478 19010
rect 14530 18958 14532 19010
rect 14476 18946 14532 18958
rect 14140 18398 14142 18450
rect 14194 18398 14196 18450
rect 14140 18386 14196 18398
rect 12012 18286 12014 18338
rect 12066 18286 12068 18338
rect 12012 18274 12068 18286
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 14812 17892 14868 19182
rect 14924 19236 14980 19246
rect 14924 18452 14980 19180
rect 15372 19236 15428 19742
rect 15484 19458 15540 20190
rect 15708 20188 15876 20244
rect 15596 20018 15652 20030
rect 15596 19966 15598 20018
rect 15650 19966 15652 20018
rect 15596 19908 15652 19966
rect 15596 19842 15652 19852
rect 15484 19406 15486 19458
rect 15538 19406 15540 19458
rect 15484 19394 15540 19406
rect 15708 19460 15764 20188
rect 15372 19170 15428 19180
rect 15708 19122 15764 19404
rect 15932 20132 15988 20142
rect 16044 20132 16100 21532
rect 16156 21586 16212 21598
rect 16156 21534 16158 21586
rect 16210 21534 16212 21586
rect 16156 21028 16212 21534
rect 16156 20804 16212 20972
rect 16156 20738 16212 20748
rect 15988 20076 16100 20132
rect 15932 20018 15988 20076
rect 15932 19966 15934 20018
rect 15986 19966 15988 20018
rect 15932 19348 15988 19966
rect 15932 19282 15988 19292
rect 15708 19070 15710 19122
rect 15762 19070 15764 19122
rect 15708 19058 15764 19070
rect 16156 19124 16212 19134
rect 15596 19012 15652 19022
rect 15596 18918 15652 18956
rect 15372 18452 15428 18462
rect 14924 18450 15428 18452
rect 14924 18398 14926 18450
rect 14978 18398 15374 18450
rect 15426 18398 15428 18450
rect 14924 18396 15428 18398
rect 14924 18386 14980 18396
rect 14812 17826 14868 17836
rect 1932 17778 1988 17790
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 16884 1988 17726
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 13468 17668 13524 17678
rect 1932 16818 1988 16828
rect 13468 16884 13524 17612
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 13468 16210 13524 16828
rect 15148 16212 15204 18396
rect 15372 18386 15428 18396
rect 16044 17892 16100 17902
rect 16044 17798 16100 17836
rect 15708 17444 15764 17454
rect 13468 16158 13470 16210
rect 13522 16158 13524 16210
rect 13468 16146 13524 16158
rect 14924 16156 15148 16212
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14924 14532 14980 16156
rect 15148 16118 15204 16156
rect 15372 17442 15764 17444
rect 15372 17390 15710 17442
rect 15762 17390 15764 17442
rect 15372 17388 15764 17390
rect 15372 17106 15428 17388
rect 15708 17378 15764 17388
rect 15372 17054 15374 17106
rect 15426 17054 15428 17106
rect 15372 15316 15428 17054
rect 16156 17106 16212 19068
rect 16268 18116 16324 25116
rect 16380 24052 16436 24062
rect 17612 24052 17668 24062
rect 16380 24050 16884 24052
rect 16380 23998 16382 24050
rect 16434 23998 16884 24050
rect 16380 23996 16884 23998
rect 16380 23986 16436 23996
rect 16828 23940 16884 23996
rect 17612 23958 17668 23996
rect 17724 23940 17780 23950
rect 16884 23884 17108 23940
rect 16828 23846 16884 23884
rect 16492 23268 16548 23278
rect 16492 22036 16548 23212
rect 17052 22372 17108 23884
rect 17164 23714 17220 23726
rect 17164 23662 17166 23714
rect 17218 23662 17220 23714
rect 17164 23156 17220 23662
rect 17724 23378 17780 23884
rect 17724 23326 17726 23378
rect 17778 23326 17780 23378
rect 17724 23314 17780 23326
rect 17836 23156 17892 26236
rect 17948 26180 18004 26460
rect 18396 26404 18452 27806
rect 18620 27188 18676 27198
rect 18732 27188 18788 27918
rect 20860 27970 20916 28364
rect 21308 28354 21364 28364
rect 20860 27918 20862 27970
rect 20914 27918 20916 27970
rect 20860 27906 20916 27918
rect 18620 27186 18788 27188
rect 18620 27134 18622 27186
rect 18674 27134 18788 27186
rect 18620 27132 18788 27134
rect 20188 27858 20244 27870
rect 20188 27806 20190 27858
rect 20242 27806 20244 27858
rect 18620 27122 18676 27132
rect 19516 27076 19572 27086
rect 18508 26404 18564 26414
rect 18396 26402 18564 26404
rect 18396 26350 18510 26402
rect 18562 26350 18564 26402
rect 18396 26348 18564 26350
rect 18508 26338 18564 26348
rect 18844 26404 18900 26414
rect 18844 26310 18900 26348
rect 18956 26402 19012 26414
rect 18956 26350 18958 26402
rect 19010 26350 19012 26402
rect 18956 26292 19012 26350
rect 18956 26226 19012 26236
rect 19180 26290 19236 26302
rect 19516 26292 19572 27020
rect 20188 26964 20244 27806
rect 20748 27188 20804 27198
rect 20188 26898 20244 26908
rect 20300 27186 20804 27188
rect 20300 27134 20750 27186
rect 20802 27134 20804 27186
rect 20300 27132 20804 27134
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20300 26516 20356 27132
rect 20748 27122 20804 27132
rect 21308 27188 21364 27198
rect 21308 27074 21364 27132
rect 21644 27186 21700 28476
rect 23996 27970 24052 27982
rect 23996 27918 23998 27970
rect 24050 27918 24052 27970
rect 23772 27858 23828 27870
rect 23772 27806 23774 27858
rect 23826 27806 23828 27858
rect 21644 27134 21646 27186
rect 21698 27134 21700 27186
rect 21644 27122 21700 27134
rect 21756 27748 21812 27758
rect 21308 27022 21310 27074
rect 21362 27022 21364 27074
rect 21308 27010 21364 27022
rect 21532 27076 21588 27086
rect 21532 26982 21588 27020
rect 21756 27074 21812 27692
rect 22988 27748 23044 27758
rect 22988 27654 23044 27692
rect 23436 27746 23492 27758
rect 23436 27694 23438 27746
rect 23490 27694 23492 27746
rect 21756 27022 21758 27074
rect 21810 27022 21812 27074
rect 21756 27010 21812 27022
rect 21980 27636 22036 27646
rect 21980 27074 22036 27580
rect 21980 27022 21982 27074
rect 22034 27022 22036 27074
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 19180 26180 19236 26238
rect 18004 26124 18340 26180
rect 17948 26114 18004 26124
rect 18172 25508 18228 25518
rect 18172 25414 18228 25452
rect 17948 25396 18004 25406
rect 17948 25302 18004 25340
rect 18284 24946 18340 26124
rect 19180 26114 19236 26124
rect 19292 26290 19572 26292
rect 19292 26238 19518 26290
rect 19570 26238 19572 26290
rect 19292 26236 19572 26238
rect 19292 25618 19348 26236
rect 19516 26226 19572 26236
rect 19964 26460 20356 26516
rect 20972 26964 21028 26974
rect 20972 26514 21028 26908
rect 20972 26462 20974 26514
rect 21026 26462 21028 26514
rect 19292 25566 19294 25618
rect 19346 25566 19348 25618
rect 19292 25554 19348 25566
rect 19068 25508 19124 25518
rect 19964 25508 20020 26460
rect 20972 26450 21028 26462
rect 21980 26514 22036 27022
rect 21980 26462 21982 26514
rect 22034 26462 22036 26514
rect 21980 26450 22036 26462
rect 22988 27076 23044 27086
rect 23436 27076 23492 27694
rect 23772 27186 23828 27806
rect 23772 27134 23774 27186
rect 23826 27134 23828 27186
rect 23772 27122 23828 27134
rect 22988 27074 23492 27076
rect 22988 27022 22990 27074
rect 23042 27022 23492 27074
rect 22988 27020 23492 27022
rect 22988 26964 23044 27020
rect 23996 26908 24052 27918
rect 24108 27860 24164 27870
rect 24108 27766 24164 27804
rect 24556 27748 24612 37998
rect 26796 37490 26852 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26796 37438 26798 37490
rect 26850 37438 26852 37490
rect 26796 37426 26852 37438
rect 25788 37266 25844 37278
rect 25788 37214 25790 37266
rect 25842 37214 25844 37266
rect 25788 31948 25844 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 25340 31892 25844 31948
rect 25340 28084 25396 31892
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 25340 28082 25956 28084
rect 25340 28030 25342 28082
rect 25394 28030 25956 28082
rect 25340 28028 25956 28030
rect 25340 28018 25396 28028
rect 25116 27860 25172 27870
rect 25116 27766 25172 27804
rect 25452 27860 25508 27870
rect 25452 27766 25508 27804
rect 24556 27682 24612 27692
rect 25900 27186 25956 28028
rect 26796 27860 26852 27870
rect 25900 27134 25902 27186
rect 25954 27134 25956 27186
rect 25900 27122 25956 27134
rect 26236 27300 26292 27310
rect 18732 25396 18788 25406
rect 18620 25284 18676 25294
rect 18620 24948 18676 25228
rect 18284 24894 18286 24946
rect 18338 24894 18340 24946
rect 18284 24882 18340 24894
rect 18508 24946 18676 24948
rect 18508 24894 18622 24946
rect 18674 24894 18676 24946
rect 18508 24892 18676 24894
rect 17164 23100 18116 23156
rect 17276 22596 17332 22606
rect 17948 22596 18004 22606
rect 17276 22594 17892 22596
rect 17276 22542 17278 22594
rect 17330 22542 17892 22594
rect 17276 22540 17892 22542
rect 17276 22530 17332 22540
rect 17164 22372 17220 22382
rect 17052 22370 17220 22372
rect 17052 22318 17166 22370
rect 17218 22318 17220 22370
rect 17052 22316 17220 22318
rect 17164 22306 17220 22316
rect 17724 22372 17780 22382
rect 16380 21812 16436 21822
rect 16380 20132 16436 21756
rect 16492 21586 16548 21980
rect 17612 22146 17668 22158
rect 17612 22094 17614 22146
rect 17666 22094 17668 22146
rect 17612 21924 17668 22094
rect 17612 21858 17668 21868
rect 17052 21700 17108 21710
rect 16492 21534 16494 21586
rect 16546 21534 16548 21586
rect 16492 21522 16548 21534
rect 16716 21588 16772 21598
rect 16492 21364 16548 21374
rect 16492 21270 16548 21308
rect 16716 20580 16772 21532
rect 16828 21364 16884 21374
rect 16828 21270 16884 21308
rect 17052 20802 17108 21644
rect 17276 21028 17332 21038
rect 17164 20972 17276 21028
rect 17164 20914 17220 20972
rect 17276 20962 17332 20972
rect 17164 20862 17166 20914
rect 17218 20862 17220 20914
rect 17164 20850 17220 20862
rect 17052 20750 17054 20802
rect 17106 20750 17108 20802
rect 17052 20738 17108 20750
rect 17276 20804 17332 20814
rect 17724 20804 17780 22316
rect 17836 21812 17892 22540
rect 17948 22502 18004 22540
rect 18060 22372 18116 23100
rect 18284 23044 18340 23054
rect 18284 23042 18452 23044
rect 18284 22990 18286 23042
rect 18338 22990 18452 23042
rect 18284 22988 18452 22990
rect 18284 22978 18340 22988
rect 18284 22372 18340 22382
rect 18060 22370 18340 22372
rect 18060 22318 18286 22370
rect 18338 22318 18340 22370
rect 18060 22316 18340 22318
rect 18284 22306 18340 22316
rect 18060 21924 18116 21934
rect 17836 21756 18004 21812
rect 17836 21586 17892 21598
rect 17836 21534 17838 21586
rect 17890 21534 17892 21586
rect 17836 21028 17892 21534
rect 17836 20962 17892 20972
rect 17724 20748 17892 20804
rect 16716 20514 16772 20524
rect 16380 20066 16436 20076
rect 16492 20468 16548 20478
rect 16268 18050 16324 18060
rect 16380 19908 16436 19918
rect 16380 18450 16436 19852
rect 16380 18398 16382 18450
rect 16434 18398 16436 18450
rect 16268 17780 16324 17790
rect 16380 17780 16436 18398
rect 16268 17778 16436 17780
rect 16268 17726 16270 17778
rect 16322 17726 16436 17778
rect 16268 17724 16436 17726
rect 16268 17714 16324 17724
rect 16492 17668 16548 20412
rect 17276 19234 17332 20748
rect 17388 20692 17444 20702
rect 17388 20598 17444 20636
rect 17724 20580 17780 20590
rect 17724 20486 17780 20524
rect 17388 20244 17444 20254
rect 17388 20132 17444 20188
rect 17500 20132 17556 20142
rect 17388 20130 17556 20132
rect 17388 20078 17502 20130
rect 17554 20078 17556 20130
rect 17388 20076 17556 20078
rect 17388 19908 17444 19918
rect 17388 19814 17444 19852
rect 17500 19572 17556 20076
rect 17724 20132 17780 20142
rect 17836 20132 17892 20748
rect 17724 20130 17892 20132
rect 17724 20078 17726 20130
rect 17778 20078 17892 20130
rect 17724 20076 17892 20078
rect 17948 20132 18004 21756
rect 18060 20802 18116 21868
rect 18060 20750 18062 20802
rect 18114 20750 18116 20802
rect 18060 20738 18116 20750
rect 18172 21698 18228 21710
rect 18172 21646 18174 21698
rect 18226 21646 18228 21698
rect 18172 21364 18228 21646
rect 18284 21700 18340 21710
rect 18396 21700 18452 22988
rect 18508 22596 18564 24892
rect 18620 24882 18676 24892
rect 18620 23268 18676 23278
rect 18732 23268 18788 25340
rect 18956 23380 19012 23390
rect 18676 23212 18788 23268
rect 18844 23324 18956 23380
rect 18620 23174 18676 23212
rect 18508 22530 18564 22540
rect 18508 22260 18564 22270
rect 18732 22260 18788 22270
rect 18508 22258 18732 22260
rect 18508 22206 18510 22258
rect 18562 22206 18732 22258
rect 18508 22204 18732 22206
rect 18508 22194 18564 22204
rect 18732 22194 18788 22204
rect 18844 22146 18900 23324
rect 18956 23286 19012 23324
rect 18844 22094 18846 22146
rect 18898 22094 18900 22146
rect 18844 21924 18900 22094
rect 18844 21858 18900 21868
rect 18956 22484 19012 22494
rect 18340 21644 18452 21700
rect 18508 21698 18564 21710
rect 18508 21646 18510 21698
rect 18562 21646 18564 21698
rect 18284 21634 18340 21644
rect 18172 20804 18228 21308
rect 18396 20804 18452 20814
rect 18172 20802 18452 20804
rect 18172 20750 18398 20802
rect 18450 20750 18452 20802
rect 18172 20748 18452 20750
rect 18172 20132 18228 20142
rect 17948 20130 18228 20132
rect 17948 20078 18174 20130
rect 18226 20078 18228 20130
rect 17948 20076 18228 20078
rect 17724 20066 17780 20076
rect 17500 19516 17892 19572
rect 17276 19182 17278 19234
rect 17330 19182 17332 19234
rect 17276 19170 17332 19182
rect 17612 19346 17668 19358
rect 17612 19294 17614 19346
rect 17666 19294 17668 19346
rect 16828 19124 16884 19134
rect 16828 19030 16884 19068
rect 17612 19124 17668 19294
rect 17612 19058 17668 19068
rect 17724 19236 17780 19246
rect 16716 18676 16772 18686
rect 16604 18562 16660 18574
rect 16604 18510 16606 18562
rect 16658 18510 16660 18562
rect 16604 18116 16660 18510
rect 16604 18050 16660 18060
rect 16156 17054 16158 17106
rect 16210 17054 16212 17106
rect 15932 16884 15988 16894
rect 15932 16790 15988 16828
rect 15484 16770 15540 16782
rect 15708 16772 15764 16782
rect 15484 16718 15486 16770
rect 15538 16718 15540 16770
rect 15484 16212 15540 16718
rect 15596 16716 15708 16772
rect 15596 16658 15652 16716
rect 15708 16706 15764 16716
rect 15596 16606 15598 16658
rect 15650 16606 15652 16658
rect 15596 16594 15652 16606
rect 15596 16212 15652 16222
rect 15484 16210 15652 16212
rect 15484 16158 15598 16210
rect 15650 16158 15652 16210
rect 15484 16156 15652 16158
rect 15596 16146 15652 16156
rect 15596 15316 15652 15326
rect 16156 15316 16212 17054
rect 16380 17612 16548 17668
rect 16380 17106 16436 17612
rect 16380 17054 16382 17106
rect 16434 17054 16436 17106
rect 16380 17042 16436 17054
rect 16492 17444 16548 17454
rect 16492 17106 16548 17388
rect 16492 17054 16494 17106
rect 16546 17054 16548 17106
rect 16492 17042 16548 17054
rect 16268 16772 16324 16782
rect 16268 16678 16324 16716
rect 16268 16212 16324 16222
rect 16268 16098 16324 16156
rect 16268 16046 16270 16098
rect 16322 16046 16324 16098
rect 16268 16034 16324 16046
rect 15372 15314 15764 15316
rect 15372 15262 15598 15314
rect 15650 15262 15764 15314
rect 15372 15260 15764 15262
rect 15596 15250 15652 15260
rect 15596 15090 15652 15102
rect 15596 15038 15598 15090
rect 15650 15038 15652 15090
rect 15596 14642 15652 15038
rect 15596 14590 15598 14642
rect 15650 14590 15652 14642
rect 15596 14578 15652 14590
rect 14028 14530 14980 14532
rect 14028 14478 14926 14530
rect 14978 14478 14980 14530
rect 14028 14476 14980 14478
rect 14028 13746 14084 14476
rect 14924 14466 14980 14476
rect 15708 14532 15764 15260
rect 15932 15204 15988 15242
rect 16156 15222 16212 15260
rect 16604 15314 16660 15326
rect 16604 15262 16606 15314
rect 16658 15262 16660 15314
rect 15932 15138 15988 15148
rect 16380 15202 16436 15214
rect 16380 15150 16382 15202
rect 16434 15150 16436 15202
rect 16380 14756 16436 15150
rect 16604 15148 16660 15262
rect 16716 15314 16772 18620
rect 17724 18562 17780 19180
rect 17836 19234 17892 19516
rect 17836 19182 17838 19234
rect 17890 19182 17892 19234
rect 17836 19170 17892 19182
rect 17724 18510 17726 18562
rect 17778 18510 17780 18562
rect 17724 18498 17780 18510
rect 17836 18452 17892 18462
rect 17948 18452 18004 20076
rect 18172 20066 18228 20076
rect 17836 18450 17948 18452
rect 17836 18398 17838 18450
rect 17890 18398 17948 18450
rect 17836 18396 17948 18398
rect 17836 18386 17892 18396
rect 17948 18358 18004 18396
rect 18060 19236 18116 19246
rect 18060 18450 18116 19180
rect 18396 19124 18452 20748
rect 18396 19058 18452 19068
rect 18508 20580 18564 21646
rect 18956 20802 19012 22428
rect 19068 21812 19124 25452
rect 19628 25506 20020 25508
rect 19628 25454 19966 25506
rect 20018 25454 20020 25506
rect 19628 25452 20020 25454
rect 19180 25396 19236 25406
rect 19180 25302 19236 25340
rect 19404 25394 19460 25406
rect 19404 25342 19406 25394
rect 19458 25342 19460 25394
rect 19292 23828 19348 23838
rect 19292 22484 19348 23772
rect 19404 23716 19460 25342
rect 19404 23650 19460 23660
rect 19516 24722 19572 24734
rect 19516 24670 19518 24722
rect 19570 24670 19572 24722
rect 19068 21698 19124 21756
rect 19068 21646 19070 21698
rect 19122 21646 19124 21698
rect 19068 21634 19124 21646
rect 19180 22482 19348 22484
rect 19180 22430 19294 22482
rect 19346 22430 19348 22482
rect 19180 22428 19348 22430
rect 19180 22260 19236 22428
rect 19292 22418 19348 22428
rect 19404 22596 19460 22606
rect 19404 22260 19460 22540
rect 18956 20750 18958 20802
rect 19010 20750 19012 20802
rect 18956 20738 19012 20750
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 18060 18386 18116 18398
rect 18284 18452 18340 18462
rect 18508 18452 18564 20524
rect 19180 20020 19236 22204
rect 19292 22204 19460 22260
rect 19292 21364 19348 22204
rect 19404 21924 19460 21934
rect 19404 21586 19460 21868
rect 19404 21534 19406 21586
rect 19458 21534 19460 21586
rect 19404 21522 19460 21534
rect 19516 21476 19572 24670
rect 19628 23380 19684 25452
rect 19964 25442 20020 25452
rect 21756 26290 21812 26302
rect 21756 26238 21758 26290
rect 21810 26238 21812 26290
rect 21756 26068 21812 26238
rect 19740 25284 19796 25322
rect 19740 25218 19796 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20636 23940 20692 23950
rect 21420 23940 21476 23950
rect 20636 23938 20804 23940
rect 20636 23886 20638 23938
rect 20690 23886 20804 23938
rect 20636 23884 20804 23886
rect 20636 23874 20692 23884
rect 20300 23828 20356 23838
rect 20300 23734 20356 23772
rect 20524 23716 20580 23726
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23324 20020 23380
rect 19292 21308 19460 21364
rect 19292 20020 19348 20030
rect 19180 19964 19292 20020
rect 19292 19954 19348 19964
rect 18620 19906 18676 19918
rect 18620 19854 18622 19906
rect 18674 19854 18676 19906
rect 18620 18676 18676 19854
rect 19404 19236 19460 21308
rect 19404 19142 19460 19180
rect 18620 18610 18676 18620
rect 19180 19124 19236 19134
rect 18956 18562 19012 18574
rect 18956 18510 18958 18562
rect 19010 18510 19012 18562
rect 18284 18450 18564 18452
rect 18284 18398 18286 18450
rect 18338 18398 18564 18450
rect 18284 18396 18564 18398
rect 18620 18452 18676 18462
rect 18284 18340 18340 18396
rect 18620 18358 18676 18396
rect 18956 18452 19012 18510
rect 18956 18386 19012 18396
rect 18284 18274 18340 18284
rect 19068 17780 19124 17790
rect 18620 17778 19124 17780
rect 18620 17726 19070 17778
rect 19122 17726 19124 17778
rect 18620 17724 19124 17726
rect 16828 16212 16884 16222
rect 16828 16118 16884 16156
rect 17836 16212 17892 16222
rect 17836 16100 17892 16156
rect 18620 16210 18676 17724
rect 19068 17714 19124 17724
rect 19180 17554 19236 19068
rect 19180 17502 19182 17554
rect 19234 17502 19236 17554
rect 19180 17490 19236 17502
rect 19292 19012 19348 19022
rect 18620 16158 18622 16210
rect 18674 16158 18676 16210
rect 18620 16146 18676 16158
rect 17612 16098 17892 16100
rect 17612 16046 17838 16098
rect 17890 16046 17892 16098
rect 17612 16044 17892 16046
rect 16716 15262 16718 15314
rect 16770 15262 16772 15314
rect 16716 15250 16772 15262
rect 17388 15316 17444 15326
rect 17388 15222 17444 15260
rect 17500 15204 17556 15242
rect 16604 15092 16772 15148
rect 17500 15138 17556 15148
rect 16716 15036 16884 15092
rect 16380 14690 16436 14700
rect 15708 14466 15764 14476
rect 14700 14308 14756 14318
rect 14700 13858 14756 14252
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13682 14084 13694
rect 16828 13634 16884 15036
rect 17612 14644 17668 16044
rect 17836 16034 17892 16044
rect 17948 15988 18004 15998
rect 17948 15426 18004 15932
rect 19292 15988 19348 18956
rect 19404 17556 19460 17566
rect 19404 17462 19460 17500
rect 19516 16882 19572 21420
rect 19628 23044 19684 23054
rect 19628 20804 19684 22988
rect 19964 23042 20020 23324
rect 19964 22990 19966 23042
rect 20018 22990 20020 23042
rect 19964 22932 20020 22990
rect 19964 22866 20020 22876
rect 20412 23042 20468 23054
rect 20412 22990 20414 23042
rect 20466 22990 20468 23042
rect 20188 22484 20244 22494
rect 20412 22484 20468 22990
rect 20188 22370 20244 22428
rect 20188 22318 20190 22370
rect 20242 22318 20244 22370
rect 20188 22306 20244 22318
rect 20300 22428 20412 22484
rect 19852 22148 19908 22186
rect 19852 22082 19908 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20300 21924 20356 22428
rect 20412 22418 20468 22428
rect 19836 21914 20100 21924
rect 20188 21868 20356 21924
rect 20076 21028 20132 21038
rect 20076 20914 20132 20972
rect 20076 20862 20078 20914
rect 20130 20862 20132 20914
rect 20076 20850 20132 20862
rect 19852 20804 19908 20814
rect 19684 20802 19908 20804
rect 19684 20750 19854 20802
rect 19906 20750 19908 20802
rect 19684 20748 19908 20750
rect 19628 20710 19684 20748
rect 19852 20738 19908 20748
rect 20076 20692 20132 20702
rect 20188 20692 20244 21868
rect 20412 21026 20468 21038
rect 20412 20974 20414 21026
rect 20466 20974 20468 21026
rect 20132 20636 20244 20692
rect 20076 20626 20132 20636
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20244 20244 20636
rect 19964 20188 20244 20244
rect 20300 20802 20356 20814
rect 20300 20750 20302 20802
rect 20354 20750 20356 20802
rect 19964 20018 20020 20188
rect 19964 19966 19966 20018
rect 20018 19966 20020 20018
rect 19964 19954 20020 19966
rect 20300 20020 20356 20750
rect 20300 19926 20356 19964
rect 19628 19346 19684 19358
rect 19628 19294 19630 19346
rect 19682 19294 19684 19346
rect 19628 18674 19684 19294
rect 19740 19122 19796 19134
rect 19740 19070 19742 19122
rect 19794 19070 19796 19122
rect 19740 19012 19796 19070
rect 19740 18946 19796 18956
rect 20300 19122 20356 19134
rect 20300 19070 20302 19122
rect 20354 19070 20356 19122
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18622 19630 18674
rect 19682 18622 19684 18674
rect 19628 18340 19684 18622
rect 19628 18274 19684 18284
rect 19964 18562 20020 18574
rect 19964 18510 19966 18562
rect 20018 18510 20020 18562
rect 19964 18228 20020 18510
rect 19964 18162 20020 18172
rect 20300 18452 20356 19070
rect 20300 17780 20356 18396
rect 19852 17724 20356 17780
rect 20412 17892 20468 20974
rect 20524 20020 20580 23660
rect 20636 23714 20692 23726
rect 20636 23662 20638 23714
rect 20690 23662 20692 23714
rect 20636 21588 20692 23662
rect 20636 21522 20692 21532
rect 20748 22370 20804 23884
rect 21420 23846 21476 23884
rect 21308 23714 21364 23726
rect 21308 23662 21310 23714
rect 21362 23662 21364 23714
rect 20860 23154 20916 23166
rect 20860 23102 20862 23154
rect 20914 23102 20916 23154
rect 20860 22932 20916 23102
rect 20860 22866 20916 22876
rect 21308 22596 21364 23662
rect 21756 23380 21812 26012
rect 22876 25620 22932 25630
rect 22316 25618 22932 25620
rect 22316 25566 22878 25618
rect 22930 25566 22932 25618
rect 22316 25564 22932 25566
rect 21868 24052 21924 24062
rect 21868 24050 22148 24052
rect 21868 23998 21870 24050
rect 21922 23998 22148 24050
rect 21868 23996 22148 23998
rect 21868 23986 21924 23996
rect 21868 23380 21924 23390
rect 21756 23378 21924 23380
rect 21756 23326 21870 23378
rect 21922 23326 21924 23378
rect 21756 23324 21924 23326
rect 21868 23314 21924 23324
rect 21756 23156 21812 23166
rect 21756 23062 21812 23100
rect 21308 22530 21364 22540
rect 21532 23042 21588 23054
rect 21532 22990 21534 23042
rect 21586 22990 21588 23042
rect 20748 22318 20750 22370
rect 20802 22318 20804 22370
rect 20748 21028 20804 22318
rect 21420 22260 21476 22270
rect 20748 20962 20804 20972
rect 21308 21924 21364 21934
rect 21308 21700 21364 21868
rect 21308 20802 21364 21644
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 21308 20738 21364 20750
rect 20524 19234 20580 19964
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 20524 19170 20580 19182
rect 20636 20132 20692 20142
rect 20636 19236 20692 20076
rect 21420 20130 21476 22204
rect 21532 21028 21588 22990
rect 22092 22260 22148 23996
rect 22316 23940 22372 25564
rect 22876 25554 22932 25564
rect 22988 24834 23044 26908
rect 23660 26852 24052 26908
rect 24668 26852 24724 26862
rect 23660 26404 23716 26852
rect 24668 26514 24724 26796
rect 24668 26462 24670 26514
rect 24722 26462 24724 26514
rect 24668 26450 24724 26462
rect 25452 26852 25508 26862
rect 23660 26310 23716 26348
rect 22988 24782 22990 24834
rect 23042 24782 23044 24834
rect 22988 24770 23044 24782
rect 23548 26290 23604 26302
rect 23548 26238 23550 26290
rect 23602 26238 23604 26290
rect 23548 24164 23604 26238
rect 23884 26292 23940 26302
rect 25452 26292 25508 26796
rect 26236 26402 26292 27244
rect 26796 26962 26852 27804
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 27468 27300 27524 27310
rect 27468 27206 27524 27244
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 26796 26910 26798 26962
rect 26850 26910 26852 26962
rect 26236 26350 26238 26402
rect 26290 26350 26292 26402
rect 26236 26338 26292 26350
rect 26348 26852 26404 26862
rect 23884 26290 25060 26292
rect 23884 26238 23886 26290
rect 23938 26238 25060 26290
rect 23884 26236 25060 26238
rect 23884 26226 23940 26236
rect 25004 25618 25060 26236
rect 25452 26290 25732 26292
rect 25452 26238 25454 26290
rect 25506 26238 25732 26290
rect 25452 26236 25732 26238
rect 25452 26226 25508 26236
rect 25004 25566 25006 25618
rect 25058 25566 25060 25618
rect 25004 25554 25060 25566
rect 25676 25508 25732 26236
rect 26236 25620 26292 25630
rect 26348 25620 26404 26796
rect 26796 26740 26852 26910
rect 26908 27076 26964 27086
rect 26908 26962 26964 27020
rect 27132 27076 27188 27086
rect 27580 27076 27636 27086
rect 27132 27074 27636 27076
rect 27132 27022 27134 27074
rect 27186 27022 27582 27074
rect 27634 27022 27636 27074
rect 27132 27020 27636 27022
rect 27132 27010 27188 27020
rect 27580 27010 27636 27020
rect 28364 27076 28420 27086
rect 26908 26910 26910 26962
rect 26962 26910 26964 26962
rect 26908 26898 26964 26910
rect 27468 26850 27524 26862
rect 27468 26798 27470 26850
rect 27522 26798 27524 26850
rect 26796 26684 26964 26740
rect 26236 25618 26404 25620
rect 26236 25566 26238 25618
rect 26290 25566 26404 25618
rect 26236 25564 26404 25566
rect 26236 25554 26292 25564
rect 25452 25506 25732 25508
rect 25452 25454 25678 25506
rect 25730 25454 25732 25506
rect 25452 25452 25732 25454
rect 26908 25508 26964 26684
rect 27020 25508 27076 25518
rect 26908 25506 27076 25508
rect 26908 25454 27022 25506
rect 27074 25454 27076 25506
rect 26908 25452 27076 25454
rect 25452 24946 25508 25452
rect 25452 24894 25454 24946
rect 25506 24894 25508 24946
rect 23660 24164 23716 24174
rect 23548 24162 23716 24164
rect 23548 24110 23662 24162
rect 23714 24110 23716 24162
rect 23548 24108 23716 24110
rect 23660 24098 23716 24108
rect 24780 24050 24836 24062
rect 24780 23998 24782 24050
rect 24834 23998 24836 24050
rect 24332 23940 24388 23950
rect 22372 23884 22820 23940
rect 22316 23846 22372 23884
rect 22764 23154 22820 23884
rect 24332 23846 24388 23884
rect 22764 23102 22766 23154
rect 22818 23102 22820 23154
rect 22764 23090 22820 23102
rect 22876 23826 22932 23838
rect 22876 23774 22878 23826
rect 22930 23774 22932 23826
rect 22876 23156 22932 23774
rect 23212 23826 23268 23838
rect 23212 23774 23214 23826
rect 23266 23774 23268 23826
rect 22988 23380 23044 23390
rect 22988 23266 23044 23324
rect 22988 23214 22990 23266
rect 23042 23214 23044 23266
rect 22988 23202 23044 23214
rect 23212 23156 23268 23774
rect 23772 23826 23828 23838
rect 23772 23774 23774 23826
rect 23826 23774 23828 23826
rect 23660 23716 23716 23726
rect 23660 23622 23716 23660
rect 23772 23268 23828 23774
rect 24780 23716 24836 23998
rect 25340 24052 25396 24062
rect 25452 24052 25508 24894
rect 25676 24724 25732 25452
rect 27020 25442 27076 25452
rect 27132 25508 27188 25518
rect 27132 25394 27188 25452
rect 27132 25342 27134 25394
rect 27186 25342 27188 25394
rect 27132 25330 27188 25342
rect 26684 25284 26740 25294
rect 25788 24724 25844 24734
rect 25676 24722 25844 24724
rect 25676 24670 25790 24722
rect 25842 24670 25844 24722
rect 25676 24668 25844 24670
rect 25788 24658 25844 24668
rect 26572 24612 26628 24622
rect 26460 24610 26628 24612
rect 26460 24558 26574 24610
rect 26626 24558 26628 24610
rect 26460 24556 26628 24558
rect 26460 24162 26516 24556
rect 26572 24546 26628 24556
rect 26460 24110 26462 24162
rect 26514 24110 26516 24162
rect 26460 24098 26516 24110
rect 25340 24050 25508 24052
rect 25340 23998 25342 24050
rect 25394 23998 25508 24050
rect 25340 23996 25508 23998
rect 25340 23986 25396 23996
rect 24780 23650 24836 23660
rect 25452 23492 25508 23996
rect 26572 23940 26628 23950
rect 26684 23940 26740 25228
rect 27356 25284 27412 25294
rect 27356 25190 27412 25228
rect 26572 23938 26740 23940
rect 26572 23886 26574 23938
rect 26626 23886 26740 23938
rect 26572 23884 26740 23886
rect 26572 23874 26628 23884
rect 26460 23716 26516 23726
rect 25340 23436 25452 23492
rect 24220 23380 24276 23390
rect 24220 23286 24276 23324
rect 23772 23202 23828 23212
rect 24108 23268 24164 23278
rect 23660 23156 23716 23166
rect 23212 23100 23660 23156
rect 22428 22930 22484 22942
rect 22428 22878 22430 22930
rect 22482 22878 22484 22930
rect 22428 22820 22484 22878
rect 22428 22754 22484 22764
rect 22876 22372 22932 23100
rect 23660 23062 23716 23100
rect 22876 22278 22932 22316
rect 23324 22930 23380 22942
rect 23324 22878 23326 22930
rect 23378 22878 23380 22930
rect 22092 22166 22148 22204
rect 23100 22258 23156 22270
rect 23100 22206 23102 22258
rect 23154 22206 23156 22258
rect 23100 21924 23156 22206
rect 23100 21858 23156 21868
rect 21868 21476 21924 21486
rect 21868 21382 21924 21420
rect 22428 21476 22484 21486
rect 21532 20934 21588 20972
rect 22316 20804 22372 20814
rect 22316 20710 22372 20748
rect 21420 20078 21422 20130
rect 21474 20078 21476 20130
rect 21420 20066 21476 20078
rect 22316 19460 22372 19470
rect 22428 19460 22484 21420
rect 22988 21026 23044 21038
rect 22988 20974 22990 21026
rect 23042 20974 23044 21026
rect 22764 20916 22820 20926
rect 22764 20130 22820 20860
rect 22876 20802 22932 20814
rect 22876 20750 22878 20802
rect 22930 20750 22932 20802
rect 22876 20244 22932 20750
rect 22988 20692 23044 20974
rect 22988 20626 23044 20636
rect 23324 20244 23380 22878
rect 23436 22932 23492 22942
rect 23436 22838 23492 22876
rect 23772 22930 23828 22942
rect 23772 22878 23774 22930
rect 23826 22878 23828 22930
rect 23772 22596 23828 22878
rect 23772 22530 23828 22540
rect 23548 22372 23604 22382
rect 23548 20802 23604 22316
rect 23548 20750 23550 20802
rect 23602 20750 23604 20802
rect 23548 20738 23604 20750
rect 23660 20916 23716 20926
rect 22876 20178 22932 20188
rect 22988 20188 23380 20244
rect 22764 20078 22766 20130
rect 22818 20078 22820 20130
rect 22764 20066 22820 20078
rect 22988 20020 23044 20188
rect 22876 20018 23044 20020
rect 22876 19966 22990 20018
rect 23042 19966 23044 20018
rect 22876 19964 23044 19966
rect 22316 19458 22708 19460
rect 22316 19406 22318 19458
rect 22370 19406 22708 19458
rect 22316 19404 22708 19406
rect 22316 19394 22372 19404
rect 20636 18674 20692 19180
rect 21980 19236 22036 19246
rect 21980 19142 22036 19180
rect 22540 19236 22596 19274
rect 22540 19170 22596 19180
rect 20636 18622 20638 18674
rect 20690 18622 20692 18674
rect 20636 18610 20692 18622
rect 21756 19124 21812 19134
rect 21756 18676 21812 19068
rect 22540 19010 22596 19022
rect 22540 18958 22542 19010
rect 22594 18958 22596 19010
rect 21756 18620 22036 18676
rect 21868 18450 21924 18462
rect 21868 18398 21870 18450
rect 21922 18398 21924 18450
rect 19740 17556 19796 17566
rect 19852 17556 19908 17724
rect 19516 16830 19518 16882
rect 19570 16830 19572 16882
rect 19516 16818 19572 16830
rect 19628 17554 19908 17556
rect 19628 17502 19742 17554
rect 19794 17502 19908 17554
rect 19628 17500 19908 17502
rect 20076 17556 20132 17566
rect 19292 15922 19348 15932
rect 17948 15374 17950 15426
rect 18002 15374 18004 15426
rect 17948 15362 18004 15374
rect 19516 15426 19572 15438
rect 19516 15374 19518 15426
rect 19570 15374 19572 15426
rect 17500 13972 17556 13982
rect 17612 13972 17668 14588
rect 17500 13970 17668 13972
rect 17500 13918 17502 13970
rect 17554 13918 17668 13970
rect 17500 13916 17668 13918
rect 17724 15314 17780 15326
rect 17724 15262 17726 15314
rect 17778 15262 17780 15314
rect 17724 14642 17780 15262
rect 19516 15316 19572 15374
rect 19628 15428 19684 17500
rect 19740 17490 19796 17500
rect 19964 17444 20020 17482
rect 20076 17462 20132 17500
rect 20300 17556 20356 17566
rect 20300 17462 20356 17500
rect 19964 17378 20020 17388
rect 20188 17442 20244 17454
rect 20188 17390 20190 17442
rect 20242 17390 20244 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 16660 20244 17390
rect 20188 16594 20244 16604
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20300 15540 20356 15550
rect 20412 15540 20468 17836
rect 20524 18228 20580 18238
rect 20524 17556 20580 18172
rect 20524 16436 20580 17500
rect 21868 17444 21924 18398
rect 21980 17556 22036 18620
rect 22540 18562 22596 18958
rect 22540 18510 22542 18562
rect 22594 18510 22596 18562
rect 22540 18498 22596 18510
rect 21980 17490 22036 17500
rect 22428 17556 22484 17566
rect 22428 17462 22484 17500
rect 21868 16994 21924 17388
rect 21868 16942 21870 16994
rect 21922 16942 21924 16994
rect 21868 16930 21924 16942
rect 20636 16660 20692 16670
rect 20692 16604 20804 16660
rect 20636 16594 20692 16604
rect 20524 16380 20692 16436
rect 20300 15538 20468 15540
rect 20300 15486 20302 15538
rect 20354 15486 20468 15538
rect 20300 15484 20468 15486
rect 20636 15538 20692 16380
rect 20748 16212 20804 16604
rect 22652 16212 22708 19404
rect 22764 17668 22820 17678
rect 22876 17668 22932 19964
rect 22988 19954 23044 19964
rect 23212 19794 23268 19806
rect 23212 19742 23214 19794
rect 23266 19742 23268 19794
rect 22764 17666 22932 17668
rect 22764 17614 22766 17666
rect 22818 17614 22932 17666
rect 22764 17612 22932 17614
rect 22988 19460 23044 19470
rect 23212 19460 23268 19742
rect 22988 19234 23044 19404
rect 22988 19182 22990 19234
rect 23042 19182 23044 19234
rect 22764 17602 22820 17612
rect 20748 16210 21364 16212
rect 20748 16158 20750 16210
rect 20802 16158 21364 16210
rect 20748 16156 21364 16158
rect 22652 16156 22932 16212
rect 20748 16146 20804 16156
rect 20636 15486 20638 15538
rect 20690 15486 20692 15538
rect 20300 15474 20356 15484
rect 20636 15474 20692 15486
rect 20076 15428 20132 15438
rect 19628 15426 20132 15428
rect 19628 15374 20078 15426
rect 20130 15374 20132 15426
rect 19628 15372 20132 15374
rect 20076 15362 20132 15372
rect 19516 15250 19572 15260
rect 20524 15314 20580 15326
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 19628 15202 19684 15214
rect 19628 15150 19630 15202
rect 19682 15150 19684 15202
rect 18060 14756 18116 14766
rect 18060 14662 18116 14700
rect 17724 14590 17726 14642
rect 17778 14590 17780 14642
rect 17500 13906 17556 13916
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16828 8428 16884 13582
rect 17724 8428 17780 14590
rect 18844 14644 18900 14654
rect 18844 14550 18900 14588
rect 19292 14644 19348 14654
rect 18396 14532 18452 14542
rect 18396 14438 18452 14476
rect 18172 14308 18228 14318
rect 18172 14214 18228 14252
rect 19292 13746 19348 14588
rect 19628 13972 19684 15150
rect 19740 15204 19796 15242
rect 19740 15138 19796 15148
rect 20412 15204 20468 15242
rect 20412 15138 20468 15148
rect 20524 15092 20580 15262
rect 21196 15314 21252 15326
rect 21196 15262 21198 15314
rect 21250 15262 21252 15314
rect 21196 15092 21252 15262
rect 20524 15036 21252 15092
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13916 20020 13972
rect 19964 13858 20020 13916
rect 19964 13806 19966 13858
rect 20018 13806 20020 13858
rect 19964 13794 20020 13806
rect 19292 13694 19294 13746
rect 19346 13694 19348 13746
rect 19292 13682 19348 13694
rect 21084 13524 21140 13534
rect 21196 13524 21252 15036
rect 21140 13468 21252 13524
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 16828 8372 17444 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 17388 4338 17444 8372
rect 17388 4286 17390 4338
rect 17442 4286 17444 4338
rect 17388 4274 17444 4286
rect 17612 8372 17780 8428
rect 16828 4116 16884 4126
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16828 800 16884 4060
rect 17500 3668 17556 3678
rect 17276 3330 17332 3342
rect 17276 3278 17278 3330
rect 17330 3278 17332 3330
rect 17276 1762 17332 3278
rect 17276 1710 17278 1762
rect 17330 1710 17332 1762
rect 17276 1698 17332 1710
rect 17500 800 17556 3612
rect 17612 3554 17668 8372
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20188 5236 20244 5246
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18396 4116 18452 4126
rect 18396 4022 18452 4060
rect 18620 3668 18676 3678
rect 18620 3574 18676 3612
rect 17612 3502 17614 3554
rect 17666 3502 17668 3554
rect 17612 3490 17668 3502
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 18172 1762 18228 1774
rect 18172 1710 18174 1762
rect 18226 1710 18228 1762
rect 18172 800 18228 1710
rect 20188 800 20244 5180
rect 21084 4338 21140 13468
rect 21308 5122 21364 16156
rect 21868 16098 21924 16110
rect 21868 16046 21870 16098
rect 21922 16046 21924 16098
rect 21532 15988 21588 15998
rect 21532 15894 21588 15932
rect 21644 15874 21700 15886
rect 21644 15822 21646 15874
rect 21698 15822 21700 15874
rect 21532 15426 21588 15438
rect 21532 15374 21534 15426
rect 21586 15374 21588 15426
rect 21532 8428 21588 15374
rect 21644 13748 21700 15822
rect 21868 15428 21924 16046
rect 21868 15362 21924 15372
rect 22316 15874 22372 15886
rect 22316 15822 22318 15874
rect 22370 15822 22372 15874
rect 21644 13682 21700 13692
rect 22316 14532 22372 15822
rect 22092 13634 22148 13646
rect 22092 13582 22094 13634
rect 22146 13582 22148 13634
rect 22092 13524 22148 13582
rect 22092 13458 22148 13468
rect 22316 13076 22372 14476
rect 22876 15316 22932 16156
rect 22988 15428 23044 19182
rect 23100 19404 23268 19460
rect 23436 19794 23492 19806
rect 23436 19742 23438 19794
rect 23490 19742 23492 19794
rect 23436 19460 23492 19742
rect 23100 19234 23156 19404
rect 23436 19394 23492 19404
rect 23548 19460 23604 19470
rect 23660 19460 23716 20860
rect 24108 20802 24164 23212
rect 25228 23268 25284 23278
rect 24444 23156 24500 23166
rect 24444 23062 24500 23100
rect 24444 22820 24500 22830
rect 24444 21028 24500 22764
rect 25228 22594 25284 23212
rect 25228 22542 25230 22594
rect 25282 22542 25284 22594
rect 24780 22484 24836 22494
rect 24836 22428 25172 22484
rect 24780 22370 24836 22428
rect 24780 22318 24782 22370
rect 24834 22318 24836 22370
rect 24780 22306 24836 22318
rect 25116 22370 25172 22428
rect 25116 22318 25118 22370
rect 25170 22318 25172 22370
rect 25116 22306 25172 22318
rect 25228 22372 25284 22542
rect 25228 22306 25284 22316
rect 24892 22260 24948 22270
rect 24892 22166 24948 22204
rect 25228 22146 25284 22158
rect 25228 22094 25230 22146
rect 25282 22094 25284 22146
rect 25228 21924 25284 22094
rect 25340 21924 25396 23436
rect 25452 23426 25508 23436
rect 26236 23714 26516 23716
rect 26236 23662 26462 23714
rect 26514 23662 26516 23714
rect 26236 23660 26516 23662
rect 25452 23156 25508 23166
rect 25452 23042 25508 23100
rect 25452 22990 25454 23042
rect 25506 22990 25508 23042
rect 25452 22978 25508 22990
rect 25676 22372 25732 22382
rect 25676 22278 25732 22316
rect 25564 22260 25620 22270
rect 25564 22036 25620 22204
rect 26236 22260 26292 23660
rect 26460 23650 26516 23660
rect 26348 23044 26404 23054
rect 26348 22594 26404 22988
rect 26348 22542 26350 22594
rect 26402 22542 26404 22594
rect 26348 22530 26404 22542
rect 26236 22166 26292 22204
rect 25788 22148 25844 22158
rect 25788 22146 25956 22148
rect 25788 22094 25790 22146
rect 25842 22094 25956 22146
rect 25788 22092 25956 22094
rect 25788 22082 25844 22092
rect 25564 21980 25732 22036
rect 25340 21868 25508 21924
rect 25228 21858 25284 21868
rect 25228 21476 25284 21486
rect 25228 21382 25284 21420
rect 24444 21026 24948 21028
rect 24444 20974 24446 21026
rect 24498 20974 24948 21026
rect 24444 20972 24948 20974
rect 24444 20962 24500 20972
rect 24220 20916 24276 20926
rect 24220 20822 24276 20860
rect 24108 20750 24110 20802
rect 24162 20750 24164 20802
rect 24108 20738 24164 20750
rect 23772 20578 23828 20590
rect 23772 20526 23774 20578
rect 23826 20526 23828 20578
rect 23772 20244 23828 20526
rect 24108 20244 24164 20254
rect 23828 20242 24164 20244
rect 23828 20190 24110 20242
rect 24162 20190 24164 20242
rect 23828 20188 24164 20190
rect 23772 20178 23828 20188
rect 24108 20178 24164 20188
rect 24444 20132 24500 20142
rect 24500 20076 24612 20132
rect 24444 20038 24500 20076
rect 23548 19458 23716 19460
rect 23548 19406 23550 19458
rect 23602 19406 23716 19458
rect 23548 19404 23716 19406
rect 23884 19794 23940 19806
rect 23884 19742 23886 19794
rect 23938 19742 23940 19794
rect 23548 19394 23604 19404
rect 23100 19182 23102 19234
rect 23154 19182 23156 19234
rect 23100 18676 23156 19182
rect 23324 19234 23380 19246
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 19124 23380 19182
rect 23324 19058 23380 19068
rect 23436 19010 23492 19022
rect 23436 18958 23438 19010
rect 23490 18958 23492 19010
rect 23436 18900 23492 18958
rect 23436 18834 23492 18844
rect 23156 18620 23604 18676
rect 23100 18610 23156 18620
rect 23324 15876 23380 15886
rect 23212 15428 23268 15438
rect 22988 15372 23212 15428
rect 23212 15334 23268 15372
rect 22876 13746 22932 15260
rect 22988 14420 23044 14430
rect 22988 14418 23268 14420
rect 22988 14366 22990 14418
rect 23042 14366 23268 14418
rect 22988 14364 23268 14366
rect 22988 14354 23044 14364
rect 23212 13970 23268 14364
rect 23212 13918 23214 13970
rect 23266 13918 23268 13970
rect 23212 13906 23268 13918
rect 22876 13694 22878 13746
rect 22930 13694 22932 13746
rect 22876 13682 22932 13694
rect 23100 13748 23156 13758
rect 23100 13654 23156 13692
rect 23324 13746 23380 15820
rect 23436 15540 23492 15550
rect 23548 15540 23604 18620
rect 23884 18452 23940 19742
rect 23884 18386 23940 18396
rect 24444 17444 24500 17454
rect 24444 17350 24500 17388
rect 24444 16324 24500 16334
rect 24556 16324 24612 20076
rect 24892 19458 24948 20972
rect 25452 20916 25508 21868
rect 25564 21698 25620 21710
rect 25564 21646 25566 21698
rect 25618 21646 25620 21698
rect 25564 21588 25620 21646
rect 25564 21522 25620 21532
rect 25676 21586 25732 21980
rect 25676 21534 25678 21586
rect 25730 21534 25732 21586
rect 25676 21522 25732 21534
rect 25788 21812 25844 21822
rect 25452 20914 25732 20916
rect 25452 20862 25454 20914
rect 25506 20862 25732 20914
rect 25452 20860 25732 20862
rect 25452 20850 25508 20860
rect 25676 20802 25732 20860
rect 25676 20750 25678 20802
rect 25730 20750 25732 20802
rect 25676 20738 25732 20750
rect 24892 19406 24894 19458
rect 24946 19406 24948 19458
rect 24892 19394 24948 19406
rect 25676 20132 25732 20142
rect 25116 19348 25172 19358
rect 25116 19254 25172 19292
rect 25452 19236 25508 19246
rect 25452 19142 25508 19180
rect 25564 19236 25620 19246
rect 25676 19236 25732 20076
rect 25788 20130 25844 21756
rect 25788 20078 25790 20130
rect 25842 20078 25844 20130
rect 25788 20066 25844 20078
rect 25564 19234 25732 19236
rect 25564 19182 25566 19234
rect 25618 19182 25732 19234
rect 25564 19180 25732 19182
rect 25564 19170 25620 19180
rect 25340 19012 25396 19022
rect 25228 18450 25284 18462
rect 25228 18398 25230 18450
rect 25282 18398 25284 18450
rect 24668 18340 24724 18350
rect 24668 18246 24724 18284
rect 25228 18116 25284 18398
rect 25340 18340 25396 18956
rect 25788 18564 25844 18574
rect 25900 18564 25956 22092
rect 26012 22146 26068 22158
rect 26012 22094 26014 22146
rect 26066 22094 26068 22146
rect 26012 22036 26068 22094
rect 26348 22146 26404 22158
rect 26348 22094 26350 22146
rect 26402 22094 26404 22146
rect 26348 22036 26404 22094
rect 26012 21980 26404 22036
rect 27468 21812 27524 26798
rect 28364 26178 28420 27020
rect 37660 27076 37716 27086
rect 37660 26982 37716 27020
rect 40012 26964 40068 27134
rect 40012 26898 40068 26908
rect 28364 26126 28366 26178
rect 28418 26126 28420 26178
rect 28364 26114 28420 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 28700 25508 28756 25518
rect 28700 24610 28756 25452
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 28700 24558 28702 24610
rect 28754 24558 28756 24610
rect 28700 24546 28756 24558
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 28252 23492 28308 23502
rect 28252 23154 28308 23436
rect 28252 23102 28254 23154
rect 28306 23102 28308 23154
rect 28252 23090 28308 23102
rect 27580 23044 27636 23054
rect 27580 22950 27636 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 27468 21746 27524 21756
rect 40236 21698 40292 21710
rect 40236 21646 40238 21698
rect 40290 21646 40292 21698
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 28588 20916 28644 20926
rect 28588 20914 29204 20916
rect 28588 20862 28590 20914
rect 28642 20862 29204 20914
rect 28588 20860 29204 20862
rect 28588 20850 28644 20860
rect 29148 20802 29204 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 29148 20750 29150 20802
rect 29202 20750 29204 20802
rect 26460 20692 26516 20702
rect 26124 20690 26516 20692
rect 26124 20638 26462 20690
rect 26514 20638 26516 20690
rect 26124 20636 26516 20638
rect 26124 20242 26180 20636
rect 26460 20626 26516 20636
rect 26124 20190 26126 20242
rect 26178 20190 26180 20242
rect 26124 20178 26180 20190
rect 27020 20132 27076 20142
rect 26012 20018 26068 20030
rect 26012 19966 26014 20018
rect 26066 19966 26068 20018
rect 26012 18900 26068 19966
rect 26236 20018 26292 20030
rect 26236 19966 26238 20018
rect 26290 19966 26292 20018
rect 26236 19796 26292 19966
rect 26460 20020 26516 20030
rect 26460 19926 26516 19964
rect 26796 20020 26852 20030
rect 26796 19926 26852 19964
rect 27020 20018 27076 20076
rect 27020 19966 27022 20018
rect 27074 19966 27076 20018
rect 27020 19954 27076 19966
rect 29148 20020 29204 20750
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 29484 20580 29540 20590
rect 29484 20486 29540 20524
rect 40012 20244 40068 20862
rect 40236 20916 40292 21646
rect 40236 20850 40292 20860
rect 40012 20178 40068 20188
rect 29148 19954 29204 19964
rect 37660 20020 37716 20030
rect 37660 19926 37716 19964
rect 26684 19906 26740 19918
rect 26684 19854 26686 19906
rect 26738 19854 26740 19906
rect 26684 19796 26740 19854
rect 26236 19740 26740 19796
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 26012 18834 26068 18844
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 26124 18564 26180 18574
rect 25900 18562 26180 18564
rect 25900 18510 26126 18562
rect 26178 18510 26180 18562
rect 25900 18508 26180 18510
rect 25788 18470 25844 18508
rect 25340 18274 25396 18284
rect 25564 18450 25620 18462
rect 25564 18398 25566 18450
rect 25618 18398 25620 18450
rect 25004 17780 25060 17790
rect 25228 17780 25284 18060
rect 25564 18116 25620 18398
rect 26012 18452 26068 18508
rect 26124 18498 26180 18508
rect 26236 18564 26292 18574
rect 26236 18470 26292 18508
rect 28252 18564 28308 18574
rect 26012 18386 26068 18396
rect 25676 18340 25732 18350
rect 25676 18338 25956 18340
rect 25676 18286 25678 18338
rect 25730 18286 25956 18338
rect 25676 18284 25956 18286
rect 25676 18274 25732 18284
rect 25564 18050 25620 18060
rect 25900 17892 25956 18284
rect 26796 18338 26852 18350
rect 26796 18286 26798 18338
rect 26850 18286 26852 18338
rect 26236 18226 26292 18238
rect 26236 18174 26238 18226
rect 26290 18174 26292 18226
rect 26236 18116 26292 18174
rect 26236 18050 26292 18060
rect 25900 17836 26180 17892
rect 25004 17778 25284 17780
rect 25004 17726 25006 17778
rect 25058 17726 25284 17778
rect 25004 17724 25284 17726
rect 26124 17778 26180 17836
rect 26124 17726 26126 17778
rect 26178 17726 26180 17778
rect 25004 17714 25060 17724
rect 26124 17714 26180 17726
rect 24444 16322 24612 16324
rect 24444 16270 24446 16322
rect 24498 16270 24612 16322
rect 24444 16268 24612 16270
rect 25340 17666 25396 17678
rect 25340 17614 25342 17666
rect 25394 17614 25396 17666
rect 25340 17444 25396 17614
rect 24220 15876 24276 15886
rect 23436 15538 23604 15540
rect 23436 15486 23438 15538
rect 23490 15486 23604 15538
rect 23436 15484 23604 15486
rect 24108 15874 24276 15876
rect 24108 15822 24222 15874
rect 24274 15822 24276 15874
rect 24108 15820 24276 15822
rect 23436 15474 23492 15484
rect 23996 15316 24052 15326
rect 23772 15314 24052 15316
rect 23772 15262 23998 15314
rect 24050 15262 24052 15314
rect 23772 15260 24052 15262
rect 23548 15204 23604 15214
rect 23772 15204 23828 15260
rect 23996 15250 24052 15260
rect 23548 15202 23828 15204
rect 23548 15150 23550 15202
rect 23602 15150 23828 15202
rect 23548 15148 23828 15150
rect 23548 15138 23604 15148
rect 23884 15090 23940 15102
rect 23884 15038 23886 15090
rect 23938 15038 23940 15090
rect 23884 14644 23940 15038
rect 24108 14756 24164 15820
rect 24220 15810 24276 15820
rect 24332 15876 24388 15886
rect 24332 15782 24388 15820
rect 24220 15316 24276 15326
rect 24220 15222 24276 15260
rect 24332 15092 24388 15102
rect 24332 14998 24388 15036
rect 24220 14756 24276 14766
rect 24108 14700 24220 14756
rect 24220 14690 24276 14700
rect 23884 14578 23940 14588
rect 23324 13694 23326 13746
rect 23378 13694 23380 13746
rect 23324 13682 23380 13694
rect 24444 13524 24500 16268
rect 25340 15540 25396 17388
rect 26796 17444 26852 18286
rect 26796 17378 26852 17388
rect 28252 17778 28308 18508
rect 37884 18450 37940 18462
rect 37884 18398 37886 18450
rect 37938 18398 37940 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 28252 17726 28254 17778
rect 28306 17726 28308 17778
rect 27916 16994 27972 17006
rect 27916 16942 27918 16994
rect 27970 16942 27972 16994
rect 27692 16884 27748 16894
rect 27692 16790 27748 16828
rect 27916 16772 27972 16942
rect 28252 16884 28308 17726
rect 28252 16818 28308 16828
rect 37660 17666 37716 17678
rect 37660 17614 37662 17666
rect 37714 17614 37716 17666
rect 27916 16706 27972 16716
rect 37660 16772 37716 17614
rect 37884 16884 37940 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 37884 16818 37940 16828
rect 37660 16706 37716 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 25788 15540 25844 15550
rect 25340 15538 25844 15540
rect 25340 15486 25342 15538
rect 25394 15486 25790 15538
rect 25842 15486 25844 15538
rect 25340 15484 25844 15486
rect 25340 15474 25396 15484
rect 25340 15092 25396 15102
rect 25116 14756 25172 14766
rect 25116 14642 25172 14700
rect 25116 14590 25118 14642
rect 25170 14590 25172 14642
rect 25116 13748 25172 14590
rect 25340 13970 25396 15036
rect 25452 14532 25508 15484
rect 25788 15474 25844 15484
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 26236 14644 26292 14654
rect 26236 14550 26292 14588
rect 28364 14642 28420 14654
rect 28364 14590 28366 14642
rect 28418 14590 28420 14642
rect 25452 14438 25508 14476
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 25340 13906 25396 13918
rect 25564 13748 25620 13758
rect 25116 13692 25396 13748
rect 24444 13458 24500 13468
rect 25228 13524 25284 13534
rect 25228 13430 25284 13468
rect 22428 13076 22484 13086
rect 22316 13074 22484 13076
rect 22316 13022 22430 13074
rect 22482 13022 22484 13074
rect 22316 13020 22484 13022
rect 22428 13010 22484 13020
rect 21308 5070 21310 5122
rect 21362 5070 21364 5122
rect 21308 5058 21364 5070
rect 21420 8372 21588 8428
rect 21084 4286 21086 4338
rect 21138 4286 21140 4338
rect 21084 4274 21140 4286
rect 20860 4116 20916 4126
rect 20860 800 20916 4060
rect 21420 3554 21476 8372
rect 22316 5236 22372 5246
rect 22316 5142 22372 5180
rect 22092 4116 22148 4126
rect 22092 4022 22148 4060
rect 21420 3502 21422 3554
rect 21474 3502 21476 3554
rect 21420 3490 21476 3502
rect 21532 3668 21588 3678
rect 21532 800 21588 3612
rect 22428 3668 22484 3678
rect 22428 3574 22484 3612
rect 24892 3668 24948 3678
rect 24892 800 24948 3612
rect 25340 3554 25396 13692
rect 25564 13654 25620 13692
rect 28364 13748 28420 14590
rect 28364 8428 28420 13692
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 27916 8372 28420 8428
rect 27916 4338 27972 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 27916 4286 27918 4338
rect 27970 4286 27972 4338
rect 27916 4274 27972 4286
rect 26012 4116 26068 4126
rect 25340 3502 25342 3554
rect 25394 3502 25396 3554
rect 25340 3490 25396 3502
rect 25564 4114 26068 4116
rect 25564 4062 26014 4114
rect 26066 4062 26068 4114
rect 25564 4060 26068 4062
rect 25564 800 25620 4060
rect 26012 4050 26068 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 26124 3668 26180 3678
rect 26124 3574 26180 3612
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 24864 0 24976 800
rect 25536 0 25648 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 25564 38556 25620 38612
rect 26796 38556 26852 38612
rect 22876 38220 22932 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 14588 28028 14644 28084
rect 4284 27858 4340 27860
rect 4284 27806 4286 27858
rect 4286 27806 4338 27858
rect 4338 27806 4340 27858
rect 4284 27804 4340 27806
rect 11788 27804 11844 27860
rect 1932 27634 1988 27636
rect 1932 27582 1934 27634
rect 1934 27582 1986 27634
rect 1986 27582 1988 27634
rect 1932 27580 1988 27582
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 1932 27186 1988 27188
rect 1932 27134 1934 27186
rect 1934 27134 1986 27186
rect 1986 27134 1988 27186
rect 1932 27132 1988 27134
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 11340 27020 11396 27076
rect 4956 26236 5012 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 1932 23548 1988 23604
rect 4284 22988 4340 23044
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 1932 21532 1988 21588
rect 15260 28082 15316 28084
rect 15260 28030 15262 28082
rect 15262 28030 15314 28082
rect 15314 28030 15316 28082
rect 15260 28028 15316 28030
rect 16940 27916 16996 27972
rect 14700 27804 14756 27860
rect 13468 25506 13524 25508
rect 13468 25454 13470 25506
rect 13470 25454 13522 25506
rect 13522 25454 13524 25506
rect 13468 25452 13524 25454
rect 14028 26348 14084 26404
rect 13692 25452 13748 25508
rect 14252 26236 14308 26292
rect 14924 26290 14980 26292
rect 14924 26238 14926 26290
rect 14926 26238 14978 26290
rect 14978 26238 14980 26290
rect 14924 26236 14980 26238
rect 15820 27804 15876 27860
rect 15372 27186 15428 27188
rect 15372 27134 15374 27186
rect 15374 27134 15426 27186
rect 15426 27134 15428 27186
rect 15372 27132 15428 27134
rect 15148 27020 15204 27076
rect 17388 27858 17444 27860
rect 17388 27806 17390 27858
rect 17390 27806 17442 27858
rect 17442 27806 17444 27858
rect 17388 27804 17444 27806
rect 16044 27020 16100 27076
rect 15372 26348 15428 26404
rect 13580 23996 13636 24052
rect 10892 23324 10948 23380
rect 14924 23996 14980 24052
rect 15260 26012 15316 26068
rect 14252 23436 14308 23492
rect 15036 23436 15092 23492
rect 14364 23378 14420 23380
rect 14364 23326 14366 23378
rect 14366 23326 14418 23378
rect 14418 23326 14420 23378
rect 14364 23324 14420 23326
rect 10892 23042 10948 23044
rect 10892 22990 10894 23042
rect 10894 22990 10946 23042
rect 10946 22990 10948 23042
rect 10892 22988 10948 22990
rect 13020 23042 13076 23044
rect 13020 22990 13022 23042
rect 13022 22990 13074 23042
rect 13074 22990 13076 23042
rect 13020 22988 13076 22990
rect 4956 22092 5012 22148
rect 14476 23154 14532 23156
rect 14476 23102 14478 23154
rect 14478 23102 14530 23154
rect 14530 23102 14532 23154
rect 14476 23100 14532 23102
rect 14364 22930 14420 22932
rect 14364 22878 14366 22930
rect 14366 22878 14418 22930
rect 14418 22878 14420 22930
rect 14364 22876 14420 22878
rect 14812 21868 14868 21924
rect 12796 21756 12852 21812
rect 14700 21810 14756 21812
rect 14700 21758 14702 21810
rect 14702 21758 14754 21810
rect 14754 21758 14756 21810
rect 14700 21756 14756 21758
rect 4284 21420 4340 21476
rect 10668 21474 10724 21476
rect 10668 21422 10670 21474
rect 10670 21422 10722 21474
rect 10722 21422 10724 21474
rect 10668 21420 10724 21422
rect 14476 21420 14532 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 15260 23436 15316 23492
rect 16044 26402 16100 26404
rect 16044 26350 16046 26402
rect 16046 26350 16098 26402
rect 16098 26350 16100 26402
rect 16044 26348 16100 26350
rect 16492 26402 16548 26404
rect 16492 26350 16494 26402
rect 16494 26350 16546 26402
rect 16546 26350 16548 26402
rect 16492 26348 16548 26350
rect 16156 25506 16212 25508
rect 16156 25454 16158 25506
rect 16158 25454 16210 25506
rect 16210 25454 16212 25506
rect 16156 25452 16212 25454
rect 15260 22988 15316 23044
rect 15148 22930 15204 22932
rect 15148 22878 15150 22930
rect 15150 22878 15202 22930
rect 15202 22878 15204 22930
rect 15148 22876 15204 22878
rect 15036 21756 15092 21812
rect 15260 21980 15316 22036
rect 14924 20860 14980 20916
rect 15260 21756 15316 21812
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 9996 19964 10052 20020
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 11676 19516 11732 19572
rect 12012 19628 12068 19684
rect 4284 19234 4340 19236
rect 4284 19182 4286 19234
rect 4286 19182 4338 19234
rect 4338 19182 4340 19234
rect 4284 19180 4340 19182
rect 14924 20578 14980 20580
rect 14924 20526 14926 20578
rect 14926 20526 14978 20578
rect 14978 20526 14980 20578
rect 14924 20524 14980 20526
rect 15148 20188 15204 20244
rect 13916 20018 13972 20020
rect 13916 19966 13918 20018
rect 13918 19966 13970 20018
rect 13970 19966 13972 20018
rect 13916 19964 13972 19966
rect 12012 19180 12068 19236
rect 1932 18844 1988 18900
rect 12908 19234 12964 19236
rect 12908 19182 12910 19234
rect 12910 19182 12962 19234
rect 12962 19182 12964 19234
rect 12908 19180 12964 19182
rect 13580 19234 13636 19236
rect 13580 19182 13582 19234
rect 13582 19182 13634 19234
rect 13634 19182 13636 19234
rect 13580 19180 13636 19182
rect 16828 26290 16884 26292
rect 16828 26238 16830 26290
rect 16830 26238 16882 26290
rect 16882 26238 16884 26290
rect 16828 26236 16884 26238
rect 16380 26124 16436 26180
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17836 28028 17892 28084
rect 17948 27970 18004 27972
rect 17948 27918 17950 27970
rect 17950 27918 18002 27970
rect 18002 27918 18004 27970
rect 17948 27916 18004 27918
rect 17724 27132 17780 27188
rect 17612 26178 17668 26180
rect 17612 26126 17614 26178
rect 17614 26126 17666 26178
rect 17666 26126 17668 26178
rect 17612 26124 17668 26126
rect 17948 26908 18004 26964
rect 17836 26290 17892 26292
rect 17836 26238 17838 26290
rect 17838 26238 17890 26290
rect 17890 26238 17892 26290
rect 17836 26236 17892 26238
rect 15708 23042 15764 23044
rect 15708 22990 15710 23042
rect 15710 22990 15762 23042
rect 15762 22990 15764 23042
rect 15708 22988 15764 22990
rect 15932 22764 15988 22820
rect 15708 21308 15764 21364
rect 15932 20802 15988 20804
rect 15932 20750 15934 20802
rect 15934 20750 15986 20802
rect 15986 20750 15988 20802
rect 15932 20748 15988 20750
rect 15708 20578 15764 20580
rect 15708 20526 15710 20578
rect 15710 20526 15762 20578
rect 15762 20526 15764 20578
rect 15708 20524 15764 20526
rect 15596 20412 15652 20468
rect 14924 19628 14980 19684
rect 14476 19516 14532 19572
rect 14140 18956 14196 19012
rect 15036 19458 15092 19460
rect 15036 19406 15038 19458
rect 15038 19406 15090 19458
rect 15090 19406 15092 19458
rect 15036 19404 15092 19406
rect 14588 19292 14644 19348
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 14924 19180 14980 19236
rect 15596 19852 15652 19908
rect 15708 19404 15764 19460
rect 15372 19180 15428 19236
rect 16156 20972 16212 21028
rect 16156 20748 16212 20804
rect 15932 20076 15988 20132
rect 15932 19292 15988 19348
rect 16156 19068 16212 19124
rect 15596 19010 15652 19012
rect 15596 18958 15598 19010
rect 15598 18958 15650 19010
rect 15650 18958 15652 19010
rect 15596 18956 15652 18958
rect 14812 17836 14868 17892
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 13468 17612 13524 17668
rect 1932 16828 1988 16884
rect 13468 16828 13524 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 16044 17890 16100 17892
rect 16044 17838 16046 17890
rect 16046 17838 16098 17890
rect 16098 17838 16100 17890
rect 16044 17836 16100 17838
rect 15148 16156 15204 16212
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 17612 24050 17668 24052
rect 17612 23998 17614 24050
rect 17614 23998 17666 24050
rect 17666 23998 17668 24050
rect 17612 23996 17668 23998
rect 16828 23938 16884 23940
rect 16828 23886 16830 23938
rect 16830 23886 16882 23938
rect 16882 23886 16884 23938
rect 16828 23884 16884 23886
rect 16492 23212 16548 23268
rect 17724 23884 17780 23940
rect 19516 27020 19572 27076
rect 18844 26402 18900 26404
rect 18844 26350 18846 26402
rect 18846 26350 18898 26402
rect 18898 26350 18900 26402
rect 18844 26348 18900 26350
rect 18956 26236 19012 26292
rect 20188 26908 20244 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 21308 27132 21364 27188
rect 21756 27692 21812 27748
rect 21532 27074 21588 27076
rect 21532 27022 21534 27074
rect 21534 27022 21586 27074
rect 21586 27022 21588 27074
rect 21532 27020 21588 27022
rect 22988 27746 23044 27748
rect 22988 27694 22990 27746
rect 22990 27694 23042 27746
rect 23042 27694 23044 27746
rect 22988 27692 23044 27694
rect 21980 27580 22036 27636
rect 17948 26124 18004 26180
rect 18172 25506 18228 25508
rect 18172 25454 18174 25506
rect 18174 25454 18226 25506
rect 18226 25454 18228 25506
rect 18172 25452 18228 25454
rect 17948 25394 18004 25396
rect 17948 25342 17950 25394
rect 17950 25342 18002 25394
rect 18002 25342 18004 25394
rect 17948 25340 18004 25342
rect 19180 26124 19236 26180
rect 20972 26908 21028 26964
rect 22988 26908 23044 26964
rect 24108 27858 24164 27860
rect 24108 27806 24110 27858
rect 24110 27806 24162 27858
rect 24162 27806 24164 27858
rect 24108 27804 24164 27806
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 25116 27858 25172 27860
rect 25116 27806 25118 27858
rect 25118 27806 25170 27858
rect 25170 27806 25172 27858
rect 25116 27804 25172 27806
rect 25452 27858 25508 27860
rect 25452 27806 25454 27858
rect 25454 27806 25506 27858
rect 25506 27806 25508 27858
rect 25452 27804 25508 27806
rect 24556 27692 24612 27748
rect 26796 27804 26852 27860
rect 26236 27244 26292 27300
rect 19068 25452 19124 25508
rect 18732 25340 18788 25396
rect 18620 25228 18676 25284
rect 17724 22370 17780 22372
rect 17724 22318 17726 22370
rect 17726 22318 17778 22370
rect 17778 22318 17780 22370
rect 17724 22316 17780 22318
rect 16492 21980 16548 22036
rect 16380 21756 16436 21812
rect 17612 21868 17668 21924
rect 17052 21644 17108 21700
rect 16716 21532 16772 21588
rect 16492 21362 16548 21364
rect 16492 21310 16494 21362
rect 16494 21310 16546 21362
rect 16546 21310 16548 21362
rect 16492 21308 16548 21310
rect 16828 21362 16884 21364
rect 16828 21310 16830 21362
rect 16830 21310 16882 21362
rect 16882 21310 16884 21362
rect 16828 21308 16884 21310
rect 17276 20972 17332 21028
rect 17276 20748 17332 20804
rect 17948 22594 18004 22596
rect 17948 22542 17950 22594
rect 17950 22542 18002 22594
rect 18002 22542 18004 22594
rect 17948 22540 18004 22542
rect 18060 21868 18116 21924
rect 17836 20972 17892 21028
rect 16716 20524 16772 20580
rect 16380 20076 16436 20132
rect 16492 20412 16548 20468
rect 16268 18060 16324 18116
rect 16380 19852 16436 19908
rect 17388 20690 17444 20692
rect 17388 20638 17390 20690
rect 17390 20638 17442 20690
rect 17442 20638 17444 20690
rect 17388 20636 17444 20638
rect 17724 20578 17780 20580
rect 17724 20526 17726 20578
rect 17726 20526 17778 20578
rect 17778 20526 17780 20578
rect 17724 20524 17780 20526
rect 17388 20188 17444 20244
rect 17388 19906 17444 19908
rect 17388 19854 17390 19906
rect 17390 19854 17442 19906
rect 17442 19854 17444 19906
rect 17388 19852 17444 19854
rect 18620 23266 18676 23268
rect 18620 23214 18622 23266
rect 18622 23214 18674 23266
rect 18674 23214 18676 23266
rect 18620 23212 18676 23214
rect 18956 23378 19012 23380
rect 18956 23326 18958 23378
rect 18958 23326 19010 23378
rect 19010 23326 19012 23378
rect 18956 23324 19012 23326
rect 18508 22540 18564 22596
rect 18732 22204 18788 22260
rect 18844 21868 18900 21924
rect 18956 22428 19012 22484
rect 18284 21644 18340 21700
rect 18172 21308 18228 21364
rect 16828 19122 16884 19124
rect 16828 19070 16830 19122
rect 16830 19070 16882 19122
rect 16882 19070 16884 19122
rect 16828 19068 16884 19070
rect 17612 19068 17668 19124
rect 17724 19180 17780 19236
rect 16716 18620 16772 18676
rect 16604 18060 16660 18116
rect 15932 16882 15988 16884
rect 15932 16830 15934 16882
rect 15934 16830 15986 16882
rect 15986 16830 15988 16882
rect 15932 16828 15988 16830
rect 15708 16716 15764 16772
rect 16492 17388 16548 17444
rect 16268 16770 16324 16772
rect 16268 16718 16270 16770
rect 16270 16718 16322 16770
rect 16322 16718 16324 16770
rect 16268 16716 16324 16718
rect 16268 16156 16324 16212
rect 16156 15314 16212 15316
rect 16156 15262 16158 15314
rect 16158 15262 16210 15314
rect 16210 15262 16212 15314
rect 16156 15260 16212 15262
rect 15932 15202 15988 15204
rect 15932 15150 15934 15202
rect 15934 15150 15986 15202
rect 15986 15150 15988 15202
rect 15932 15148 15988 15150
rect 17948 18396 18004 18452
rect 18060 19180 18116 19236
rect 18396 19068 18452 19124
rect 19180 25394 19236 25396
rect 19180 25342 19182 25394
rect 19182 25342 19234 25394
rect 19234 25342 19236 25394
rect 19180 25340 19236 25342
rect 19292 23772 19348 23828
rect 19404 23660 19460 23716
rect 19068 21756 19124 21812
rect 19404 22540 19460 22596
rect 19180 22204 19236 22260
rect 18508 20524 18564 20580
rect 19404 21868 19460 21924
rect 21756 26012 21812 26068
rect 19740 25282 19796 25284
rect 19740 25230 19742 25282
rect 19742 25230 19794 25282
rect 19794 25230 19796 25282
rect 19740 25228 19796 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 23826 20356 23828
rect 20300 23774 20302 23826
rect 20302 23774 20354 23826
rect 20354 23774 20356 23826
rect 20300 23772 20356 23774
rect 20524 23660 20580 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19516 21420 19572 21476
rect 19292 19964 19348 20020
rect 19404 19234 19460 19236
rect 19404 19182 19406 19234
rect 19406 19182 19458 19234
rect 19458 19182 19460 19234
rect 19404 19180 19460 19182
rect 18620 18620 18676 18676
rect 19180 19068 19236 19124
rect 18620 18450 18676 18452
rect 18620 18398 18622 18450
rect 18622 18398 18674 18450
rect 18674 18398 18676 18450
rect 18620 18396 18676 18398
rect 18956 18396 19012 18452
rect 18284 18284 18340 18340
rect 16828 16210 16884 16212
rect 16828 16158 16830 16210
rect 16830 16158 16882 16210
rect 16882 16158 16884 16210
rect 16828 16156 16884 16158
rect 17836 16156 17892 16212
rect 19292 18956 19348 19012
rect 17388 15314 17444 15316
rect 17388 15262 17390 15314
rect 17390 15262 17442 15314
rect 17442 15262 17444 15314
rect 17388 15260 17444 15262
rect 17500 15202 17556 15204
rect 17500 15150 17502 15202
rect 17502 15150 17554 15202
rect 17554 15150 17556 15202
rect 17500 15148 17556 15150
rect 16380 14700 16436 14756
rect 15708 14476 15764 14532
rect 14700 14252 14756 14308
rect 17948 15932 18004 15988
rect 19404 17554 19460 17556
rect 19404 17502 19406 17554
rect 19406 17502 19458 17554
rect 19458 17502 19460 17554
rect 19404 17500 19460 17502
rect 19628 23042 19684 23044
rect 19628 22990 19630 23042
rect 19630 22990 19682 23042
rect 19682 22990 19684 23042
rect 19628 22988 19684 22990
rect 19964 22876 20020 22932
rect 20188 22428 20244 22484
rect 20412 22428 20468 22484
rect 19852 22146 19908 22148
rect 19852 22094 19854 22146
rect 19854 22094 19906 22146
rect 19906 22094 19908 22146
rect 19852 22092 19908 22094
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 20972 20132 21028
rect 19628 20748 19684 20804
rect 20076 20636 20132 20692
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20300 20018 20356 20020
rect 20300 19966 20302 20018
rect 20302 19966 20354 20018
rect 20354 19966 20356 20018
rect 20300 19964 20356 19966
rect 19740 18956 19796 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18284 19684 18340
rect 19964 18172 20020 18228
rect 20300 18450 20356 18452
rect 20300 18398 20302 18450
rect 20302 18398 20354 18450
rect 20354 18398 20356 18450
rect 20300 18396 20356 18398
rect 20636 21532 20692 21588
rect 21420 23938 21476 23940
rect 21420 23886 21422 23938
rect 21422 23886 21474 23938
rect 21474 23886 21476 23938
rect 21420 23884 21476 23886
rect 20860 22876 20916 22932
rect 21756 23154 21812 23156
rect 21756 23102 21758 23154
rect 21758 23102 21810 23154
rect 21810 23102 21812 23154
rect 21756 23100 21812 23102
rect 21308 22540 21364 22596
rect 21420 22204 21476 22260
rect 20748 20972 20804 21028
rect 21308 21868 21364 21924
rect 21308 21644 21364 21700
rect 20524 19964 20580 20020
rect 20636 20076 20692 20132
rect 24668 26796 24724 26852
rect 25452 26796 25508 26852
rect 23660 26402 23716 26404
rect 23660 26350 23662 26402
rect 23662 26350 23714 26402
rect 23714 26350 23716 26402
rect 23660 26348 23716 26350
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 27468 27298 27524 27300
rect 27468 27246 27470 27298
rect 27470 27246 27522 27298
rect 27522 27246 27524 27298
rect 27468 27244 27524 27246
rect 26348 26850 26404 26852
rect 26348 26798 26350 26850
rect 26350 26798 26402 26850
rect 26402 26798 26404 26850
rect 26348 26796 26404 26798
rect 26908 27020 26964 27076
rect 28364 27020 28420 27076
rect 22316 23938 22372 23940
rect 22316 23886 22318 23938
rect 22318 23886 22370 23938
rect 22370 23886 22372 23938
rect 22316 23884 22372 23886
rect 24332 23938 24388 23940
rect 24332 23886 24334 23938
rect 24334 23886 24386 23938
rect 24386 23886 24388 23938
rect 24332 23884 24388 23886
rect 22988 23324 23044 23380
rect 22876 23100 22932 23156
rect 23660 23714 23716 23716
rect 23660 23662 23662 23714
rect 23662 23662 23714 23714
rect 23714 23662 23716 23714
rect 23660 23660 23716 23662
rect 27132 25452 27188 25508
rect 26684 25228 26740 25284
rect 24780 23660 24836 23716
rect 27356 25282 27412 25284
rect 27356 25230 27358 25282
rect 27358 25230 27410 25282
rect 27410 25230 27412 25282
rect 27356 25228 27412 25230
rect 25452 23436 25508 23492
rect 24220 23378 24276 23380
rect 24220 23326 24222 23378
rect 24222 23326 24274 23378
rect 24274 23326 24276 23378
rect 24220 23324 24276 23326
rect 23772 23212 23828 23268
rect 24108 23212 24164 23268
rect 23660 23154 23716 23156
rect 23660 23102 23662 23154
rect 23662 23102 23714 23154
rect 23714 23102 23716 23154
rect 23660 23100 23716 23102
rect 22428 22764 22484 22820
rect 22876 22370 22932 22372
rect 22876 22318 22878 22370
rect 22878 22318 22930 22370
rect 22930 22318 22932 22370
rect 22876 22316 22932 22318
rect 22092 22258 22148 22260
rect 22092 22206 22094 22258
rect 22094 22206 22146 22258
rect 22146 22206 22148 22258
rect 22092 22204 22148 22206
rect 23100 21868 23156 21924
rect 21868 21474 21924 21476
rect 21868 21422 21870 21474
rect 21870 21422 21922 21474
rect 21922 21422 21924 21474
rect 21868 21420 21924 21422
rect 22428 21420 22484 21476
rect 21532 21026 21588 21028
rect 21532 20974 21534 21026
rect 21534 20974 21586 21026
rect 21586 20974 21588 21026
rect 21532 20972 21588 20974
rect 22316 20802 22372 20804
rect 22316 20750 22318 20802
rect 22318 20750 22370 20802
rect 22370 20750 22372 20802
rect 22316 20748 22372 20750
rect 22764 20860 22820 20916
rect 22988 20636 23044 20692
rect 23436 22930 23492 22932
rect 23436 22878 23438 22930
rect 23438 22878 23490 22930
rect 23490 22878 23492 22930
rect 23436 22876 23492 22878
rect 23772 22540 23828 22596
rect 23548 22316 23604 22372
rect 23660 20860 23716 20916
rect 22876 20188 22932 20244
rect 20636 19180 20692 19236
rect 21980 19234 22036 19236
rect 21980 19182 21982 19234
rect 21982 19182 22034 19234
rect 22034 19182 22036 19234
rect 21980 19180 22036 19182
rect 22540 19234 22596 19236
rect 22540 19182 22542 19234
rect 22542 19182 22594 19234
rect 22594 19182 22596 19234
rect 22540 19180 22596 19182
rect 21756 19122 21812 19124
rect 21756 19070 21758 19122
rect 21758 19070 21810 19122
rect 21810 19070 21812 19122
rect 21756 19068 21812 19070
rect 20412 17836 20468 17892
rect 20076 17554 20132 17556
rect 20076 17502 20078 17554
rect 20078 17502 20130 17554
rect 20130 17502 20132 17554
rect 20076 17500 20132 17502
rect 19292 15932 19348 15988
rect 17612 14588 17668 14644
rect 20300 17554 20356 17556
rect 20300 17502 20302 17554
rect 20302 17502 20354 17554
rect 20354 17502 20356 17554
rect 20300 17500 20356 17502
rect 19964 17442 20020 17444
rect 19964 17390 19966 17442
rect 19966 17390 20018 17442
rect 20018 17390 20020 17442
rect 19964 17388 20020 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20188 16604 20244 16660
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20524 18172 20580 18228
rect 20524 17500 20580 17556
rect 21980 17500 22036 17556
rect 22428 17554 22484 17556
rect 22428 17502 22430 17554
rect 22430 17502 22482 17554
rect 22482 17502 22484 17554
rect 22428 17500 22484 17502
rect 21868 17388 21924 17444
rect 20636 16604 20692 16660
rect 22988 19404 23044 19460
rect 19516 15260 19572 15316
rect 18060 14754 18116 14756
rect 18060 14702 18062 14754
rect 18062 14702 18114 14754
rect 18114 14702 18116 14754
rect 18060 14700 18116 14702
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 18844 14642 18900 14644
rect 18844 14590 18846 14642
rect 18846 14590 18898 14642
rect 18898 14590 18900 14642
rect 18844 14588 18900 14590
rect 19292 14588 19348 14644
rect 18396 14530 18452 14532
rect 18396 14478 18398 14530
rect 18398 14478 18450 14530
rect 18450 14478 18452 14530
rect 18396 14476 18452 14478
rect 18172 14306 18228 14308
rect 18172 14254 18174 14306
rect 18174 14254 18226 14306
rect 18226 14254 18228 14306
rect 18172 14252 18228 14254
rect 19740 15202 19796 15204
rect 19740 15150 19742 15202
rect 19742 15150 19794 15202
rect 19794 15150 19796 15202
rect 19740 15148 19796 15150
rect 20412 15202 20468 15204
rect 20412 15150 20414 15202
rect 20414 15150 20466 15202
rect 20466 15150 20468 15202
rect 20412 15148 20468 15150
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21084 13468 21140 13524
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 16828 4060 16884 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 17500 3612 17556 3668
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20188 5180 20244 5236
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18396 4114 18452 4116
rect 18396 4062 18398 4114
rect 18398 4062 18450 4114
rect 18450 4062 18452 4114
rect 18396 4060 18452 4062
rect 18620 3666 18676 3668
rect 18620 3614 18622 3666
rect 18622 3614 18674 3666
rect 18674 3614 18676 3666
rect 18620 3612 18676 3614
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21532 15986 21588 15988
rect 21532 15934 21534 15986
rect 21534 15934 21586 15986
rect 21586 15934 21588 15986
rect 21532 15932 21588 15934
rect 21868 15372 21924 15428
rect 21644 13692 21700 13748
rect 22316 14530 22372 14532
rect 22316 14478 22318 14530
rect 22318 14478 22370 14530
rect 22370 14478 22372 14530
rect 22316 14476 22372 14478
rect 22092 13468 22148 13524
rect 23436 19404 23492 19460
rect 25228 23212 25284 23268
rect 24444 23154 24500 23156
rect 24444 23102 24446 23154
rect 24446 23102 24498 23154
rect 24498 23102 24500 23154
rect 24444 23100 24500 23102
rect 24444 22764 24500 22820
rect 24780 22428 24836 22484
rect 25228 22316 25284 22372
rect 24892 22258 24948 22260
rect 24892 22206 24894 22258
rect 24894 22206 24946 22258
rect 24946 22206 24948 22258
rect 24892 22204 24948 22206
rect 25228 21868 25284 21924
rect 25452 23100 25508 23156
rect 25676 22370 25732 22372
rect 25676 22318 25678 22370
rect 25678 22318 25730 22370
rect 25730 22318 25732 22370
rect 25676 22316 25732 22318
rect 25564 22204 25620 22260
rect 26348 22988 26404 23044
rect 26236 22258 26292 22260
rect 26236 22206 26238 22258
rect 26238 22206 26290 22258
rect 26290 22206 26292 22258
rect 26236 22204 26292 22206
rect 25228 21474 25284 21476
rect 25228 21422 25230 21474
rect 25230 21422 25282 21474
rect 25282 21422 25284 21474
rect 25228 21420 25284 21422
rect 24220 20914 24276 20916
rect 24220 20862 24222 20914
rect 24222 20862 24274 20914
rect 24274 20862 24276 20914
rect 24220 20860 24276 20862
rect 23772 20188 23828 20244
rect 24444 20130 24500 20132
rect 24444 20078 24446 20130
rect 24446 20078 24498 20130
rect 24498 20078 24500 20130
rect 24444 20076 24500 20078
rect 23324 19068 23380 19124
rect 23436 18844 23492 18900
rect 23100 18620 23156 18676
rect 23324 15820 23380 15876
rect 23212 15426 23268 15428
rect 23212 15374 23214 15426
rect 23214 15374 23266 15426
rect 23266 15374 23268 15426
rect 23212 15372 23268 15374
rect 22876 15260 22932 15316
rect 23100 13746 23156 13748
rect 23100 13694 23102 13746
rect 23102 13694 23154 13746
rect 23154 13694 23156 13746
rect 23100 13692 23156 13694
rect 23884 18396 23940 18452
rect 24444 17442 24500 17444
rect 24444 17390 24446 17442
rect 24446 17390 24498 17442
rect 24498 17390 24500 17442
rect 24444 17388 24500 17390
rect 25564 21532 25620 21588
rect 25788 21756 25844 21812
rect 25676 20076 25732 20132
rect 25116 19346 25172 19348
rect 25116 19294 25118 19346
rect 25118 19294 25170 19346
rect 25170 19294 25172 19346
rect 25116 19292 25172 19294
rect 25452 19234 25508 19236
rect 25452 19182 25454 19234
rect 25454 19182 25506 19234
rect 25506 19182 25508 19234
rect 25452 19180 25508 19182
rect 25340 19010 25396 19012
rect 25340 18958 25342 19010
rect 25342 18958 25394 19010
rect 25394 18958 25396 19010
rect 25340 18956 25396 18958
rect 24668 18338 24724 18340
rect 24668 18286 24670 18338
rect 24670 18286 24722 18338
rect 24722 18286 24724 18338
rect 24668 18284 24724 18286
rect 25788 18562 25844 18564
rect 25788 18510 25790 18562
rect 25790 18510 25842 18562
rect 25842 18510 25844 18562
rect 25788 18508 25844 18510
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 40012 26908 40068 26964
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 28700 25452 28756 25508
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 40012 24892 40068 24948
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 28252 23436 28308 23492
rect 27580 23042 27636 23044
rect 27580 22990 27582 23042
rect 27582 22990 27634 23042
rect 27634 22990 27636 23042
rect 27580 22988 27636 22990
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 27468 21756 27524 21812
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 27020 20076 27076 20132
rect 26460 20018 26516 20020
rect 26460 19966 26462 20018
rect 26462 19966 26514 20018
rect 26514 19966 26516 20018
rect 26460 19964 26516 19966
rect 26796 20018 26852 20020
rect 26796 19966 26798 20018
rect 26798 19966 26850 20018
rect 26850 19966 26852 20018
rect 26796 19964 26852 19966
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 29484 20578 29540 20580
rect 29484 20526 29486 20578
rect 29486 20526 29538 20578
rect 29538 20526 29540 20578
rect 29484 20524 29540 20526
rect 40236 20860 40292 20916
rect 40012 20188 40068 20244
rect 29148 19964 29204 20020
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 26012 18844 26068 18900
rect 40012 18844 40068 18900
rect 25340 18284 25396 18340
rect 25228 18060 25284 18116
rect 26236 18562 26292 18564
rect 26236 18510 26238 18562
rect 26238 18510 26290 18562
rect 26290 18510 26292 18562
rect 26236 18508 26292 18510
rect 28252 18508 28308 18564
rect 26012 18396 26068 18452
rect 25564 18060 25620 18116
rect 26236 18060 26292 18116
rect 25340 17388 25396 17444
rect 24332 15874 24388 15876
rect 24332 15822 24334 15874
rect 24334 15822 24386 15874
rect 24386 15822 24388 15874
rect 24332 15820 24388 15822
rect 24220 15314 24276 15316
rect 24220 15262 24222 15314
rect 24222 15262 24274 15314
rect 24274 15262 24276 15314
rect 24220 15260 24276 15262
rect 24332 15090 24388 15092
rect 24332 15038 24334 15090
rect 24334 15038 24386 15090
rect 24386 15038 24388 15090
rect 24332 15036 24388 15038
rect 24220 14700 24276 14756
rect 23884 14588 23940 14644
rect 26796 17388 26852 17444
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 27692 16882 27748 16884
rect 27692 16830 27694 16882
rect 27694 16830 27746 16882
rect 27746 16830 27748 16882
rect 27692 16828 27748 16830
rect 28252 16828 28308 16884
rect 27916 16716 27972 16772
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 40012 17500 40068 17556
rect 37884 16828 37940 16884
rect 37660 16716 37716 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 25340 15036 25396 15092
rect 25116 14700 25172 14756
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 26236 14642 26292 14644
rect 26236 14590 26238 14642
rect 26238 14590 26290 14642
rect 26290 14590 26292 14642
rect 26236 14588 26292 14590
rect 25452 14530 25508 14532
rect 25452 14478 25454 14530
rect 25454 14478 25506 14530
rect 25506 14478 25508 14530
rect 25452 14476 25508 14478
rect 24444 13468 24500 13524
rect 25228 13522 25284 13524
rect 25228 13470 25230 13522
rect 25230 13470 25282 13522
rect 25282 13470 25284 13522
rect 25228 13468 25284 13470
rect 20860 4060 20916 4116
rect 22316 5234 22372 5236
rect 22316 5182 22318 5234
rect 22318 5182 22370 5234
rect 22370 5182 22372 5234
rect 22316 5180 22372 5182
rect 22092 4114 22148 4116
rect 22092 4062 22094 4114
rect 22094 4062 22146 4114
rect 22146 4062 22148 4114
rect 22092 4060 22148 4062
rect 21532 3612 21588 3668
rect 22428 3666 22484 3668
rect 22428 3614 22430 3666
rect 22430 3614 22482 3666
rect 22482 3614 22484 3666
rect 22428 3612 22484 3614
rect 24892 3612 24948 3668
rect 25564 13746 25620 13748
rect 25564 13694 25566 13746
rect 25566 13694 25618 13746
rect 25618 13694 25620 13746
rect 25564 13692 25620 13694
rect 28364 13692 28420 13748
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 26124 3666 26180 3668
rect 26124 3614 26126 3666
rect 26126 3614 26178 3666
rect 26178 3614 26180 3666
rect 26124 3612 26180 3614
<< metal3 >>
rect 25554 38556 25564 38612
rect 25620 38556 26796 38612
rect 26852 38556 26862 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 14578 28028 14588 28084
rect 14644 28028 15260 28084
rect 15316 28028 17836 28084
rect 17892 28028 17902 28084
rect 16930 27916 16940 27972
rect 16996 27916 17948 27972
rect 18004 27916 18014 27972
rect 4274 27804 4284 27860
rect 4340 27804 11788 27860
rect 11844 27804 14700 27860
rect 14756 27804 14766 27860
rect 15810 27804 15820 27860
rect 15876 27804 17388 27860
rect 17444 27804 17454 27860
rect 24098 27804 24108 27860
rect 24164 27804 25116 27860
rect 25172 27804 25182 27860
rect 25442 27804 25452 27860
rect 25508 27804 26796 27860
rect 26852 27804 26862 27860
rect 21746 27692 21756 27748
rect 21812 27692 22988 27748
rect 23044 27692 24556 27748
rect 24612 27692 24622 27748
rect 0 27636 800 27664
rect 25452 27636 25508 27804
rect 0 27580 1932 27636
rect 1988 27580 1998 27636
rect 21970 27580 21980 27636
rect 22036 27580 25508 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 26226 27244 26236 27300
rect 26292 27244 27468 27300
rect 27524 27244 27534 27300
rect 1922 27132 1932 27188
rect 1988 27132 1998 27188
rect 15362 27132 15372 27188
rect 15428 27132 17724 27188
rect 17780 27132 17790 27188
rect 17948 27132 21308 27188
rect 21364 27132 21374 27188
rect 0 26964 800 26992
rect 1932 26964 1988 27132
rect 17948 27076 18004 27132
rect 4274 27020 4284 27076
rect 4340 27020 11340 27076
rect 11396 27020 15148 27076
rect 15204 27020 15214 27076
rect 16034 27020 16044 27076
rect 16100 27020 18004 27076
rect 19506 27020 19516 27076
rect 19572 27020 21532 27076
rect 21588 27020 21598 27076
rect 26898 27020 26908 27076
rect 26964 27020 28364 27076
rect 28420 27020 37660 27076
rect 37716 27020 37726 27076
rect 41200 26964 42000 26992
rect 0 26908 1988 26964
rect 17938 26908 17948 26964
rect 18004 26908 20188 26964
rect 20244 26908 20972 26964
rect 21028 26908 22988 26964
rect 23044 26908 23492 26964
rect 40002 26908 40012 26964
rect 40068 26908 42000 26964
rect 0 26880 800 26908
rect 23436 26852 23492 26908
rect 41200 26880 42000 26908
rect 23436 26796 24668 26852
rect 24724 26796 25452 26852
rect 25508 26796 26348 26852
rect 26404 26796 26414 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 14018 26348 14028 26404
rect 14084 26348 15372 26404
rect 15428 26348 16044 26404
rect 16100 26348 16492 26404
rect 16548 26348 16558 26404
rect 18834 26348 18844 26404
rect 18900 26348 23660 26404
rect 23716 26348 23726 26404
rect 0 26292 800 26320
rect 0 26236 4956 26292
rect 5012 26236 5022 26292
rect 14242 26236 14252 26292
rect 14308 26236 14924 26292
rect 14980 26236 14990 26292
rect 16818 26236 16828 26292
rect 16884 26236 17836 26292
rect 17892 26236 18956 26292
rect 19012 26236 19022 26292
rect 0 26208 800 26236
rect 16370 26124 16380 26180
rect 16436 26124 17612 26180
rect 17668 26124 17948 26180
rect 18004 26124 19180 26180
rect 19236 26124 19246 26180
rect 15250 26012 15260 26068
rect 15316 26012 21756 26068
rect 21812 26012 21822 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 13458 25452 13468 25508
rect 13524 25452 13692 25508
rect 13748 25452 16156 25508
rect 16212 25452 16222 25508
rect 18162 25452 18172 25508
rect 18228 25452 19068 25508
rect 19124 25452 19134 25508
rect 27122 25452 27132 25508
rect 27188 25452 28700 25508
rect 28756 25452 37660 25508
rect 37716 25452 37726 25508
rect 17938 25340 17948 25396
rect 18004 25340 18732 25396
rect 18788 25340 19180 25396
rect 19236 25340 19246 25396
rect 18610 25228 18620 25284
rect 18676 25228 19740 25284
rect 19796 25228 19806 25284
rect 26674 25228 26684 25284
rect 26740 25228 27356 25284
rect 27412 25228 27422 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 41200 24948 42000 24976
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 41200 24864 42000 24892
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 13570 23996 13580 24052
rect 13636 23996 14924 24052
rect 14980 23996 17612 24052
rect 17668 23996 17678 24052
rect 16818 23884 16828 23940
rect 16884 23884 17724 23940
rect 17780 23884 17790 23940
rect 21410 23884 21420 23940
rect 21476 23884 22316 23940
rect 22372 23884 24332 23940
rect 24388 23884 24398 23940
rect 19282 23772 19292 23828
rect 19348 23772 20300 23828
rect 20356 23772 20366 23828
rect 19394 23660 19404 23716
rect 19460 23660 20524 23716
rect 20580 23660 23660 23716
rect 23716 23660 24780 23716
rect 24836 23660 24846 23716
rect 0 23604 800 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 14242 23436 14252 23492
rect 14308 23436 15036 23492
rect 15092 23436 15102 23492
rect 15250 23436 15260 23492
rect 15316 23436 15326 23492
rect 25442 23436 25452 23492
rect 25508 23436 28252 23492
rect 28308 23436 28318 23492
rect 10882 23324 10892 23380
rect 10948 23324 14364 23380
rect 14420 23324 14430 23380
rect 15260 23156 15316 23436
rect 18946 23324 18956 23380
rect 19012 23324 22988 23380
rect 23044 23324 24220 23380
rect 24276 23324 24286 23380
rect 16482 23212 16492 23268
rect 16548 23212 18620 23268
rect 18676 23212 18686 23268
rect 23762 23212 23772 23268
rect 23828 23212 24108 23268
rect 24164 23212 25228 23268
rect 25284 23212 25294 23268
rect 14466 23100 14476 23156
rect 14532 23100 15316 23156
rect 21746 23100 21756 23156
rect 21812 23100 22876 23156
rect 22932 23100 22942 23156
rect 23650 23100 23660 23156
rect 23716 23100 24444 23156
rect 24500 23100 25452 23156
rect 25508 23100 25518 23156
rect 4274 22988 4284 23044
rect 4340 22988 10892 23044
rect 10948 22988 10958 23044
rect 13010 22988 13020 23044
rect 13076 22988 15260 23044
rect 15316 22988 15326 23044
rect 15698 22988 15708 23044
rect 15764 22988 19628 23044
rect 19684 22988 19694 23044
rect 26338 22988 26348 23044
rect 26404 22988 27580 23044
rect 27636 22988 27646 23044
rect 14354 22876 14364 22932
rect 14420 22876 15148 22932
rect 15204 22876 15214 22932
rect 19954 22876 19964 22932
rect 20020 22876 20860 22932
rect 20916 22876 23436 22932
rect 23492 22876 23502 22932
rect 15922 22764 15932 22820
rect 15988 22764 22428 22820
rect 22484 22764 24444 22820
rect 24500 22764 24510 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 17938 22540 17948 22596
rect 18004 22540 18508 22596
rect 18564 22540 19404 22596
rect 19460 22540 19470 22596
rect 20188 22540 21308 22596
rect 21364 22540 23772 22596
rect 23828 22540 23838 22596
rect 20188 22484 20244 22540
rect 18946 22428 18956 22484
rect 19012 22428 20188 22484
rect 20244 22428 20254 22484
rect 20402 22428 20412 22484
rect 20468 22428 24780 22484
rect 24836 22428 24846 22484
rect 17714 22316 17724 22372
rect 17780 22316 21476 22372
rect 22866 22316 22876 22372
rect 22932 22316 23548 22372
rect 23604 22316 23614 22372
rect 25218 22316 25228 22372
rect 25284 22316 25676 22372
rect 25732 22316 25742 22372
rect 21420 22260 21476 22316
rect 18722 22204 18732 22260
rect 18788 22204 19180 22260
rect 19236 22204 19246 22260
rect 21410 22204 21420 22260
rect 21476 22204 22092 22260
rect 22148 22204 22158 22260
rect 24882 22204 24892 22260
rect 24948 22204 25564 22260
rect 25620 22204 26236 22260
rect 26292 22204 26302 22260
rect 4946 22092 4956 22148
rect 5012 22092 19852 22148
rect 19908 22092 19918 22148
rect 15250 21980 15260 22036
rect 15316 21980 16492 22036
rect 16548 21980 16558 22036
rect 19404 21924 19460 22092
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 14802 21868 14812 21924
rect 14868 21868 17612 21924
rect 17668 21868 17678 21924
rect 18050 21868 18060 21924
rect 18116 21868 18844 21924
rect 18900 21868 18910 21924
rect 19394 21868 19404 21924
rect 19460 21868 19470 21924
rect 21298 21868 21308 21924
rect 21364 21868 23100 21924
rect 23156 21868 25228 21924
rect 25284 21868 25294 21924
rect 12786 21756 12796 21812
rect 12852 21756 14700 21812
rect 14756 21756 14766 21812
rect 15026 21756 15036 21812
rect 15092 21756 15260 21812
rect 15316 21756 16380 21812
rect 16436 21756 16446 21812
rect 19058 21756 19068 21812
rect 19124 21756 25788 21812
rect 25844 21756 27468 21812
rect 27524 21756 27534 21812
rect 17042 21644 17052 21700
rect 17108 21644 18284 21700
rect 18340 21644 21308 21700
rect 21364 21644 21374 21700
rect 0 21588 800 21616
rect 0 21532 1932 21588
rect 1988 21532 1998 21588
rect 16706 21532 16716 21588
rect 16772 21532 20636 21588
rect 20692 21532 25564 21588
rect 25620 21532 25630 21588
rect 0 21504 800 21532
rect 4274 21420 4284 21476
rect 4340 21420 10668 21476
rect 10724 21420 14476 21476
rect 14532 21420 14542 21476
rect 19506 21420 19516 21476
rect 19572 21420 21868 21476
rect 21924 21420 21934 21476
rect 22418 21420 22428 21476
rect 22484 21420 25228 21476
rect 25284 21420 25294 21476
rect 15698 21308 15708 21364
rect 15764 21308 16492 21364
rect 16548 21308 16558 21364
rect 16818 21308 16828 21364
rect 16884 21308 18172 21364
rect 18228 21308 18238 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 16146 20972 16156 21028
rect 16212 20972 17276 21028
rect 17332 20972 17836 21028
rect 17892 20972 17902 21028
rect 20066 20972 20076 21028
rect 20132 20972 20748 21028
rect 20804 20972 21532 21028
rect 21588 20972 21598 21028
rect 41200 20916 42000 20944
rect 14914 20860 14924 20916
rect 14980 20860 22764 20916
rect 22820 20860 23660 20916
rect 23716 20860 24220 20916
rect 24276 20860 24286 20916
rect 40226 20860 40236 20916
rect 40292 20860 42000 20916
rect 41200 20832 42000 20860
rect 15922 20748 15932 20804
rect 15988 20748 16156 20804
rect 16212 20748 16222 20804
rect 17266 20748 17276 20804
rect 17332 20748 19628 20804
rect 19684 20748 22316 20804
rect 22372 20748 22382 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 17378 20636 17388 20692
rect 17444 20636 20076 20692
rect 20132 20636 20142 20692
rect 22950 20636 22988 20692
rect 23044 20636 23054 20692
rect 31892 20580 31948 20748
rect 14914 20524 14924 20580
rect 14980 20524 15708 20580
rect 15764 20524 16716 20580
rect 16772 20524 16782 20580
rect 17714 20524 17724 20580
rect 17780 20524 18508 20580
rect 18564 20524 18574 20580
rect 29474 20524 29484 20580
rect 29540 20524 31948 20580
rect 15586 20412 15596 20468
rect 15652 20412 16492 20468
rect 16548 20412 16558 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 41200 20244 42000 20272
rect 15138 20188 15148 20244
rect 15204 20188 15214 20244
rect 17378 20188 17388 20244
rect 17444 20188 22876 20244
rect 22932 20188 23772 20244
rect 23828 20188 23838 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 15148 20132 15204 20188
rect 41200 20160 42000 20188
rect 15148 20076 15932 20132
rect 15988 20076 15998 20132
rect 16370 20076 16380 20132
rect 16436 20076 20636 20132
rect 20692 20076 20702 20132
rect 24434 20076 24444 20132
rect 24500 20076 25676 20132
rect 25732 20076 27020 20132
rect 27076 20076 27086 20132
rect 4274 19964 4284 20020
rect 4340 19964 9996 20020
rect 10052 19964 13916 20020
rect 13972 19964 13982 20020
rect 19282 19964 19292 20020
rect 19348 19964 20300 20020
rect 20356 19964 20366 20020
rect 20514 19964 20524 20020
rect 20580 19964 26460 20020
rect 26516 19964 26526 20020
rect 26786 19964 26796 20020
rect 26852 19964 29148 20020
rect 29204 19964 37660 20020
rect 37716 19964 37726 20020
rect 15586 19852 15596 19908
rect 15652 19852 16380 19908
rect 16436 19852 17388 19908
rect 17444 19852 17454 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 12002 19628 12012 19684
rect 12068 19628 14924 19684
rect 14980 19628 14990 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 0 19516 1988 19572
rect 11666 19516 11676 19572
rect 11732 19516 14476 19572
rect 14532 19516 14542 19572
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 0 19488 800 19516
rect 41200 19488 42000 19516
rect 15026 19404 15036 19460
rect 15092 19404 15708 19460
rect 15764 19404 15774 19460
rect 22950 19404 22988 19460
rect 23044 19404 23436 19460
rect 23492 19404 23502 19460
rect 14578 19292 14588 19348
rect 14644 19292 15148 19348
rect 15922 19292 15932 19348
rect 15988 19292 25116 19348
rect 25172 19292 25182 19348
rect 15092 19236 15148 19292
rect 4274 19180 4284 19236
rect 4340 19180 12012 19236
rect 12068 19180 12078 19236
rect 12898 19180 12908 19236
rect 12964 19180 13580 19236
rect 13636 19180 14924 19236
rect 14980 19180 14990 19236
rect 15092 19180 15372 19236
rect 15428 19180 17724 19236
rect 17780 19180 17790 19236
rect 18050 19180 18060 19236
rect 18116 19180 19404 19236
rect 19460 19180 19470 19236
rect 20626 19180 20636 19236
rect 20692 19180 21980 19236
rect 22036 19180 22046 19236
rect 22530 19180 22540 19236
rect 22596 19180 25452 19236
rect 25508 19180 25518 19236
rect 31892 19180 37660 19236
rect 37716 19180 37726 19236
rect 16146 19068 16156 19124
rect 16212 19068 16828 19124
rect 16884 19068 16894 19124
rect 17602 19068 17612 19124
rect 17668 19068 18396 19124
rect 18452 19068 19180 19124
rect 19236 19068 19246 19124
rect 21746 19068 21756 19124
rect 21812 19068 23324 19124
rect 23380 19068 23390 19124
rect 31892 19012 31948 19180
rect 14130 18956 14140 19012
rect 14196 18956 15596 19012
rect 15652 18956 15662 19012
rect 19282 18956 19292 19012
rect 19348 18956 19740 19012
rect 19796 18956 19806 19012
rect 25330 18956 25340 19012
rect 25396 18956 31948 19012
rect 0 18900 800 18928
rect 41200 18900 42000 18928
rect 0 18844 1932 18900
rect 1988 18844 1998 18900
rect 23426 18844 23436 18900
rect 23492 18844 26012 18900
rect 26068 18844 26078 18900
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 16706 18620 16716 18676
rect 16772 18620 18620 18676
rect 18676 18620 23100 18676
rect 23156 18620 23166 18676
rect 25778 18508 25788 18564
rect 25844 18508 25854 18564
rect 26226 18508 26236 18564
rect 26292 18508 28252 18564
rect 28308 18508 28318 18564
rect 25788 18452 25844 18508
rect 17938 18396 17948 18452
rect 18004 18396 18620 18452
rect 18676 18396 18686 18452
rect 18946 18396 18956 18452
rect 19012 18396 20300 18452
rect 20356 18396 20366 18452
rect 23874 18396 23884 18452
rect 23940 18396 25844 18452
rect 26002 18396 26012 18452
rect 26068 18396 26078 18452
rect 18274 18284 18284 18340
rect 18340 18284 19628 18340
rect 19684 18284 19694 18340
rect 24658 18284 24668 18340
rect 24724 18284 25340 18340
rect 25396 18284 25406 18340
rect 26012 18228 26068 18396
rect 41200 18228 42000 18256
rect 19954 18172 19964 18228
rect 20020 18172 20524 18228
rect 20580 18172 26068 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 16258 18060 16268 18116
rect 16324 18060 16604 18116
rect 16660 18060 25228 18116
rect 25284 18060 25294 18116
rect 25554 18060 25564 18116
rect 25620 18060 26236 18116
rect 26292 18060 26302 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 14802 17836 14812 17892
rect 14868 17836 16044 17892
rect 16100 17836 20412 17892
rect 20468 17836 20478 17892
rect 4274 17612 4284 17668
rect 4340 17612 13468 17668
rect 13524 17612 13534 17668
rect 41200 17556 42000 17584
rect 19394 17500 19404 17556
rect 19460 17500 20076 17556
rect 20132 17500 20142 17556
rect 20290 17500 20300 17556
rect 20356 17500 20524 17556
rect 20580 17500 20590 17556
rect 21196 17500 21980 17556
rect 22036 17500 22428 17556
rect 22484 17500 22494 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 21196 17444 21252 17500
rect 41200 17472 42000 17500
rect 16482 17388 16492 17444
rect 16548 17388 19964 17444
rect 20020 17388 21252 17444
rect 21858 17388 21868 17444
rect 21924 17388 24444 17444
rect 24500 17388 25340 17444
rect 25396 17388 26796 17444
rect 26852 17388 26862 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 0 16884 800 16912
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 13458 16828 13468 16884
rect 13524 16828 15932 16884
rect 15988 16828 15998 16884
rect 27682 16828 27692 16884
rect 27748 16828 28252 16884
rect 28308 16828 37884 16884
rect 37940 16828 37950 16884
rect 0 16800 800 16828
rect 15698 16716 15708 16772
rect 15764 16716 16268 16772
rect 16324 16716 16334 16772
rect 27906 16716 27916 16772
rect 27972 16716 37660 16772
rect 37716 16716 37726 16772
rect 20178 16604 20188 16660
rect 20244 16604 20636 16660
rect 20692 16604 20702 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 15138 16156 15148 16212
rect 15204 16156 16268 16212
rect 16324 16156 16828 16212
rect 16884 16156 17836 16212
rect 17892 16156 17902 16212
rect 17938 15932 17948 15988
rect 18004 15932 19292 15988
rect 19348 15932 21532 15988
rect 21588 15932 21598 15988
rect 23314 15820 23324 15876
rect 23380 15820 24332 15876
rect 24388 15820 24398 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 21858 15372 21868 15428
rect 21924 15372 23212 15428
rect 23268 15372 23278 15428
rect 16146 15260 16156 15316
rect 16212 15260 17388 15316
rect 17444 15260 17454 15316
rect 19506 15260 19516 15316
rect 19572 15260 22876 15316
rect 22932 15260 24220 15316
rect 24276 15260 24286 15316
rect 15922 15148 15932 15204
rect 15988 15148 17500 15204
rect 17556 15148 17566 15204
rect 19730 15148 19740 15204
rect 19796 15148 20412 15204
rect 20468 15148 20478 15204
rect 24322 15036 24332 15092
rect 24388 15036 25340 15092
rect 25396 15036 25406 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 16370 14700 16380 14756
rect 16436 14700 18060 14756
rect 18116 14700 18126 14756
rect 24210 14700 24220 14756
rect 24276 14700 25116 14756
rect 25172 14700 25182 14756
rect 17602 14588 17612 14644
rect 17668 14588 18844 14644
rect 18900 14588 19292 14644
rect 19348 14588 20188 14644
rect 23874 14588 23884 14644
rect 23940 14588 26236 14644
rect 26292 14588 26302 14644
rect 20132 14532 20188 14588
rect 15698 14476 15708 14532
rect 15764 14476 18396 14532
rect 18452 14476 18462 14532
rect 20132 14476 22316 14532
rect 22372 14476 25452 14532
rect 25508 14476 25518 14532
rect 14690 14252 14700 14308
rect 14756 14252 18172 14308
rect 18228 14252 18238 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 21634 13692 21644 13748
rect 21700 13692 23100 13748
rect 23156 13692 23166 13748
rect 25554 13692 25564 13748
rect 25620 13692 28364 13748
rect 28420 13692 28430 13748
rect 21074 13468 21084 13524
rect 21140 13468 22092 13524
rect 22148 13468 22158 13524
rect 24434 13468 24444 13524
rect 24500 13468 25228 13524
rect 25284 13468 25294 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 20178 5180 20188 5236
rect 20244 5180 22316 5236
rect 22372 5180 22382 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 16818 4060 16828 4116
rect 16884 4060 18396 4116
rect 18452 4060 18462 4116
rect 20850 4060 20860 4116
rect 20916 4060 22092 4116
rect 22148 4060 22158 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 17490 3612 17500 3668
rect 17556 3612 18620 3668
rect 18676 3612 18686 3668
rect 21522 3612 21532 3668
rect 21588 3612 22428 3668
rect 22484 3612 22494 3668
rect 24882 3612 24892 3668
rect 24948 3612 26124 3668
rect 26180 3612 26190 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 22988 20636 23044 20692
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 22988 19404 23044 19460
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 22988 20692 23044 20702
rect 22988 19460 23044 20636
rect 22988 19394 23044 19404
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24752 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18256 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21616 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _109_
timestamp 1698175906
transform 1 0 17584 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21056 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17584 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23408 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _114_
timestamp 1698175906
transform 1 0 20048 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22176 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform 1 0 21504 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26656 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_
timestamp 1698175906
transform -1 0 27776 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17024 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 18480 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 16688 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 20272 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 18816 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1698175906
transform 1 0 18256 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform -1 0 19152 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _128_
timestamp 1698175906
transform 1 0 24192 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698175906
transform -1 0 19600 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19600 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_
timestamp 1698175906
transform 1 0 24976 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform -1 0 23968 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform 1 0 23408 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 19488 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform 1 0 25536 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _136_
timestamp 1698175906
transform -1 0 22512 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform 1 0 26096 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24080 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 22960 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19600 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _142_
timestamp 1698175906
transform -1 0 19600 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform 1 0 23296 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform -1 0 17920 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _146_
timestamp 1698175906
transform -1 0 18368 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 17024 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 16352 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _149_
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform -1 0 25648 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform -1 0 24304 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _152_
timestamp 1698175906
transform -1 0 20160 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23184 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 14672 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _156_
timestamp 1698175906
transform 1 0 18704 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20720 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _158_
timestamp 1698175906
transform -1 0 16464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18368 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22176 0 -1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform 1 0 17920 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _163_
timestamp 1698175906
transform -1 0 16352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _164_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _165_
timestamp 1698175906
transform -1 0 21616 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform 1 0 25984 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _167_
timestamp 1698175906
transform -1 0 24640 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23296 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22624 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _170_
timestamp 1698175906
transform -1 0 25984 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _171_
timestamp 1698175906
transform 1 0 23072 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19936 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _173_
timestamp 1698175906
transform -1 0 26096 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _174_
timestamp 1698175906
transform 1 0 23968 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _175_
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _176_
timestamp 1698175906
transform -1 0 24640 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _177_
timestamp 1698175906
transform 1 0 19936 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _178_
timestamp 1698175906
transform -1 0 19936 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24752 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21616 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20720 0 1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _182_
timestamp 1698175906
transform 1 0 21392 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform -1 0 24640 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _184_
timestamp 1698175906
transform -1 0 23520 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _185_
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _186_
timestamp 1698175906
transform -1 0 16128 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _187_
timestamp 1698175906
transform 1 0 15792 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1698175906
transform -1 0 15792 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform -1 0 16688 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform -1 0 15008 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13552 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 15456 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _193_
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _194_
timestamp 1698175906
transform -1 0 16128 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _195_
timestamp 1698175906
transform -1 0 18480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16016 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _198_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22736 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _199_
timestamp 1698175906
transform 1 0 26432 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _200_
timestamp 1698175906
transform -1 0 26432 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _201_
timestamp 1698175906
transform -1 0 18704 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _202_
timestamp 1698175906
transform -1 0 14448 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _203_
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _204_
timestamp 1698175906
transform 1 0 11424 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _205_
timestamp 1698175906
transform -1 0 17024 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _206_
timestamp 1698175906
transform 1 0 14336 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _207_
timestamp 1698175906
transform -1 0 15680 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1698175906
transform 1 0 26880 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform -1 0 26768 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 17696 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 25984 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform -1 0 28560 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 17696 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 14448 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 14000 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 19936 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 25200 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 25312 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 19040 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 21616 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 14672 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 16576 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform -1 0 14896 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform -1 0 14448 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform -1 0 15120 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 25536 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform -1 0 13776 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 25648 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _237_
timestamp 1698175906
transform 1 0 27440 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _238_
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _239_
timestamp 1698175906
transform 1 0 21056 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__A2
timestamp 1698175906
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__B
timestamp 1698175906
transform -1 0 25088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__A2
timestamp 1698175906
transform 1 0 16912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 17584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 26208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 25312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 22288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform -1 0 17920 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 26320 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 14000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 23408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 24416 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform -1 0 22512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 26768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 25760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 18816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 14896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 15232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 15344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform -1 0 25536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 14000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 25424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 19824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 18816 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 19264 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_168
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_172
timestamp 1698175906
transform 1 0 20608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_174
timestamp 1698175906
transform 1 0 20832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_201 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23856 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 28560 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_203
timestamp 1698175906
transform 1 0 24080 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_235
timestamp 1698175906
transform 1 0 27664 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698175906
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698175906
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_189
timestamp 1698175906
transform 1 0 22512 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_221 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26096 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_237
timestamp 1698175906
transform 1 0 27888 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_146
timestamp 1698175906
transform 1 0 17696 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_154
timestamp 1698175906
transform 1 0 18592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_187
timestamp 1698175906
transform 1 0 22288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_189
timestamp 1698175906
transform 1 0 22512 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_198
timestamp 1698175906
transform 1 0 23520 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_218
timestamp 1698175906
transform 1 0 25760 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_250
timestamp 1698175906
transform 1 0 29344 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_266
timestamp 1698175906
transform 1 0 31136 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698175906
transform 1 0 32032 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698175906
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_154
timestamp 1698175906
transform 1 0 18592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_158
timestamp 1698175906
transform 1 0 19040 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1698175906
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_150
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1698175906
transform 1 0 19040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_175
timestamp 1698175906
transform 1 0 20944 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_182
timestamp 1698175906
transform 1 0 21728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_190
timestamp 1698175906
transform 1 0 22624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698175906
transform 1 0 25536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_220
timestamp 1698175906
transform 1 0 25984 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_252
timestamp 1698175906
transform 1 0 29568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_268
timestamp 1698175906
transform 1 0 31360 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_140
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_144
timestamp 1698175906
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_189
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_197
timestamp 1698175906
transform 1 0 23408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_201
timestamp 1698175906
transform 1 0 23856 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_208
timestamp 1698175906
transform 1 0 24640 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698175906
transform 1 0 28224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_120
timestamp 1698175906
transform 1 0 14784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_122
timestamp 1698175906
transform 1 0 15008 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_154
timestamp 1698175906
transform 1 0 18592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_228
timestamp 1698175906
transform 1 0 26880 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_232
timestamp 1698175906
transform 1 0 27328 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_239
timestamp 1698175906
transform 1 0 28112 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_271
timestamp 1698175906
transform 1 0 31696 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698175906
transform 1 0 15120 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_135
timestamp 1698175906
transform 1 0 16464 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_151
timestamp 1698175906
transform 1 0 18256 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_155
timestamp 1698175906
transform 1 0 18704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1698175906
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_193
timestamp 1698175906
transform 1 0 22960 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_201
timestamp 1698175906
transform 1 0 23856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_205
timestamp 1698175906
transform 1 0 24304 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_208
timestamp 1698175906
transform 1 0 24640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_212
timestamp 1698175906
transform 1 0 25088 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698175906
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_92
timestamp 1698175906
transform 1 0 11648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_123
timestamp 1698175906
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_127
timestamp 1698175906
transform 1 0 15568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_131
timestamp 1698175906
transform 1 0 16016 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_159
timestamp 1698175906
transform 1 0 19152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_161
timestamp 1698175906
transform 1 0 19376 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_174
timestamp 1698175906
transform 1 0 20832 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_178
timestamp 1698175906
transform 1 0 21280 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_180
timestamp 1698175906
transform 1 0 21504 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_225
timestamp 1698175906
transform 1 0 26544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_229
timestamp 1698175906
transform 1 0 26992 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_261
timestamp 1698175906
transform 1 0 30576 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 9520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_131
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_135
timestamp 1698175906
transform 1 0 16464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_152
timestamp 1698175906
transform 1 0 18368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_201
timestamp 1698175906
transform 1 0 23856 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_219
timestamp 1698175906
transform 1 0 25872 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_235
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_96
timestamp 1698175906
transform 1 0 12096 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_108
timestamp 1698175906
transform 1 0 13440 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_110
timestamp 1698175906
transform 1 0 13664 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_117
timestamp 1698175906
transform 1 0 14448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_119
timestamp 1698175906
transform 1 0 14672 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_131
timestamp 1698175906
transform 1 0 16016 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_148
timestamp 1698175906
transform 1 0 17920 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_186
timestamp 1698175906
transform 1 0 22176 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_232
timestamp 1698175906
transform 1 0 27328 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_264
timestamp 1698175906
transform 1 0 30912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_132
timestamp 1698175906
transform 1 0 16128 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_136
timestamp 1698175906
transform 1 0 16576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_138
timestamp 1698175906
transform 1 0 16800 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_208
timestamp 1698175906
transform 1 0 24640 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_212
timestamp 1698175906
transform 1 0 25088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_253
timestamp 1698175906
transform 1 0 29680 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_285
timestamp 1698175906
transform 1 0 33264 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_301
timestamp 1698175906
transform 1 0 35056 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698175906
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698175906
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_111
timestamp 1698175906
transform 1 0 13776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_115
timestamp 1698175906
transform 1 0 14224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_117
timestamp 1698175906
transform 1 0 14448 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_159
timestamp 1698175906
transform 1 0 19152 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_221
timestamp 1698175906
transform 1 0 26096 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_253
timestamp 1698175906
transform 1 0 29680 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_269
timestamp 1698175906
transform 1 0 31472 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_330
timestamp 1698175906
transform 1 0 38304 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_338
timestamp 1698175906
transform 1 0 39200 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_342
timestamp 1698175906
transform 1 0 39648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_344
timestamp 1698175906
transform 1 0 39872 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_131
timestamp 1698175906
transform 1 0 16016 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_139
timestamp 1698175906
transform 1 0 16912 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_163
timestamp 1698175906
transform 1 0 19600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_226
timestamp 1698175906
transform 1 0 26656 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_113
timestamp 1698175906
transform 1 0 14000 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_119
timestamp 1698175906
transform 1 0 14672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_121
timestamp 1698175906
transform 1 0 14896 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698175906
transform 1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698175906
transform 1 0 17472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_159
timestamp 1698175906
transform 1 0 19152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_161
timestamp 1698175906
transform 1 0 19376 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_186
timestamp 1698175906
transform 1 0 22176 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_243
timestamp 1698175906
transform 1 0 28560 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_275
timestamp 1698175906
transform 1 0 32144 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_136
timestamp 1698175906
transform 1 0 16576 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_143
timestamp 1698175906
transform 1 0 17360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_147
timestamp 1698175906
transform 1 0 17808 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_163
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_165
timestamp 1698175906
transform 1 0 19824 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_189
timestamp 1698175906
transform 1 0 22512 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_202
timestamp 1698175906
transform 1 0 23968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_212
timestamp 1698175906
transform 1 0 25088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_216
timestamp 1698175906
transform 1 0 25536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_220
timestamp 1698175906
transform 1 0 25984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_227
timestamp 1698175906
transform 1 0 26768 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_214
timestamp 1698175906
transform 1 0 25312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_246
timestamp 1698175906
transform 1 0 28896 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_115
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_119
timestamp 1698175906
transform 1 0 14672 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_123
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_131
timestamp 1698175906
transform 1 0 16016 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_137
timestamp 1698175906
transform 1 0 16688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_141
timestamp 1698175906
transform 1 0 17136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_152
timestamp 1698175906
transform 1 0 18368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_156
timestamp 1698175906
transform 1 0 18816 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_169
timestamp 1698175906
transform 1 0 20272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698175906
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_189
timestamp 1698175906
transform 1 0 22512 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_220
timestamp 1698175906
transform 1 0 25984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_224
timestamp 1698175906
transform 1 0 26432 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_233
timestamp 1698175906
transform 1 0 27440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_126
timestamp 1698175906
transform 1 0 15456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_128
timestamp 1698175906
transform 1 0 15680 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_155
timestamp 1698175906
transform 1 0 18704 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_163
timestamp 1698175906
transform 1 0 19600 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_177
timestamp 1698175906
transform 1 0 21168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_179
timestamp 1698175906
transform 1 0 21392 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_186
timestamp 1698175906
transform 1 0 22176 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_194
timestamp 1698175906
transform 1 0 23072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_196
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_202
timestamp 1698175906
transform 1 0 23968 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_206
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_243
timestamp 1698175906
transform 1 0 28560 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_275
timestamp 1698175906
transform 1 0 32144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_186
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_190
timestamp 1698175906
transform 1 0 22624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_221
timestamp 1698175906
transform 1 0 26096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_225
timestamp 1698175906
transform 1 0 26544 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_236
timestamp 1698175906
transform 1 0 27776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_28
timestamp 1698175906
transform 1 0 4480 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_60
timestamp 1698175906
transform 1 0 8064 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698175906
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_122
timestamp 1698175906
transform 1 0 15008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_126
timestamp 1698175906
transform 1 0 15456 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_134
timestamp 1698175906
transform 1 0 16352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_157
timestamp 1698175906
transform 1 0 18928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_165
timestamp 1698175906
transform 1 0 19824 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_195
timestamp 1698175906
transform 1 0 23184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_199
timestamp 1698175906
transform 1 0 23632 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_205
timestamp 1698175906
transform 1 0 24304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_217
timestamp 1698175906
transform 1 0 25648 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_249
timestamp 1698175906
transform 1 0 29232 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_265
timestamp 1698175906
transform 1 0 31024 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_273
timestamp 1698175906
transform 1 0 31920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_277
timestamp 1698175906
transform 1 0 32368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_139
timestamp 1698175906
transform 1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_143
timestamp 1698175906
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_145
timestamp 1698175906
transform 1 0 17584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_148
timestamp 1698175906
transform 1 0 17920 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_164
timestamp 1698175906
transform 1 0 19712 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_181
timestamp 1698175906
transform 1 0 21616 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698175906
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 32144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita58_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita58_26
timestamp 1698175906
transform 1 0 17024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 24976 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 28560 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 20944 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 25536 41200 25648 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal3 25088 14616 25088 14616 0 _000_
rlabel metal2 19992 13888 19992 13888 0 _001_
rlabel metal2 22568 18760 22568 18760 0 _002_
rlabel metal2 23240 14168 23240 14168 0 _003_
rlabel metal2 15624 14840 15624 14840 0 _004_
rlabel metal2 15568 16184 15568 16184 0 _005_
rlabel metal2 13832 26600 13832 26600 0 _006_
rlabel metal2 13552 27720 13552 27720 0 _007_
rlabel metal2 14168 18704 14168 18704 0 _008_
rlabel metal2 26152 20440 26152 20440 0 _009_
rlabel metal2 12152 19712 12152 19712 0 _010_
rlabel metal2 12824 21728 12824 21728 0 _011_
rlabel metal2 26488 24360 26488 24360 0 _012_
rlabel metal3 26880 27272 26880 27272 0 _013_
rlabel metal2 15288 21728 15288 21728 0 _014_
rlabel metal2 18704 27160 18704 27160 0 _015_
rlabel metal2 25032 25928 25032 25928 0 _016_
rlabel metal2 26376 22792 26376 22792 0 _017_
rlabel metal2 18648 16968 18648 16968 0 _018_
rlabel metal3 16576 27160 16576 27160 0 _019_
rlabel metal2 23800 27496 23800 27496 0 _020_
rlabel metal2 15288 22960 15288 22960 0 _021_
rlabel metal2 14728 14056 14728 14056 0 _022_
rlabel metal2 20888 28168 20888 28168 0 _023_
rlabel metal2 26152 17808 26152 17808 0 _024_
rlabel metal3 14784 22904 14784 22904 0 _025_
rlabel metal2 20328 20384 20328 20384 0 _026_
rlabel metal2 20384 15512 20384 15512 0 _027_
rlabel metal3 17080 14504 17080 14504 0 _028_
rlabel metal2 16184 18088 16184 18088 0 _029_
rlabel metal2 23576 17080 23576 17080 0 _030_
rlabel metal3 17248 14728 17248 14728 0 _031_
rlabel metal2 21336 27104 21336 27104 0 _032_
rlabel metal2 21672 27832 21672 27832 0 _033_
rlabel metal2 25592 18256 25592 18256 0 _034_
rlabel metal2 22792 20496 22792 20496 0 _035_
rlabel metal2 21896 15736 21896 15736 0 _036_
rlabel metal3 25816 18480 25816 18480 0 _037_
rlabel metal2 23912 15288 23912 15288 0 _038_
rlabel metal2 20664 22624 20664 22624 0 _039_
rlabel metal2 22400 19432 22400 19432 0 _040_
rlabel metal3 24864 13496 24864 13496 0 _041_
rlabel metal2 25368 14504 25368 14504 0 _042_
rlabel metal3 20104 15176 20104 15176 0 _043_
rlabel metal3 24024 19208 24024 19208 0 _044_
rlabel metal3 19768 15960 19768 15960 0 _045_
rlabel metal3 22400 13720 22400 13720 0 _046_
rlabel metal3 23856 15848 23856 15848 0 _047_
rlabel metal3 16744 15176 16744 15176 0 _048_
rlabel metal2 15624 16688 15624 16688 0 _049_
rlabel metal2 13720 26152 13720 26152 0 _050_
rlabel metal2 14448 27048 14448 27048 0 _051_
rlabel metal2 14168 25872 14168 25872 0 _052_
rlabel metal2 15736 19656 15736 19656 0 _053_
rlabel metal2 15400 19488 15400 19488 0 _054_
rlabel metal2 15512 19824 15512 19824 0 _055_
rlabel metal2 23464 18928 23464 18928 0 _056_
rlabel metal2 26264 19880 26264 19880 0 _057_
rlabel metal2 17640 22008 17640 22008 0 _058_
rlabel metal2 14280 19208 14280 19208 0 _059_
rlabel metal2 11704 19768 11704 19768 0 _060_
rlabel metal2 15512 21448 15512 21448 0 _061_
rlabel metal2 15064 21112 15064 21112 0 _062_
rlabel metal2 26712 24584 26712 24584 0 _063_
rlabel metal2 23016 23296 23016 23296 0 _064_
rlabel metal2 19656 18984 19656 18984 0 _065_
rlabel metal2 20216 22400 20216 22400 0 _066_
rlabel metal2 17640 19208 17640 19208 0 _067_
rlabel metal2 18368 23016 18368 23016 0 _068_
rlabel metal2 24808 22400 24808 22400 0 _069_
rlabel metal2 17192 20944 17192 20944 0 _070_
rlabel metal2 27496 24304 27496 24304 0 _071_
rlabel metal3 23240 22344 23240 22344 0 _072_
rlabel metal2 20104 20944 20104 20944 0 _073_
rlabel metal2 14952 27832 14952 27832 0 _074_
rlabel metal2 26936 26096 26936 26096 0 _075_
rlabel metal2 27384 27048 27384 27048 0 _076_
rlabel metal2 18088 20104 18088 20104 0 _077_
rlabel metal2 19712 17528 19712 17528 0 _078_
rlabel metal2 17192 23408 17192 23408 0 _079_
rlabel metal2 18648 25088 18648 25088 0 _080_
rlabel metal3 17024 26152 17024 26152 0 _081_
rlabel metal2 18480 26376 18480 26376 0 _082_
rlabel metal2 16520 21784 16520 21784 0 _083_
rlabel metal3 21560 23688 21560 23688 0 _084_
rlabel metal3 20552 27048 20552 27048 0 _085_
rlabel metal2 24024 27412 24024 27412 0 _086_
rlabel metal2 25256 22904 25256 22904 0 _087_
rlabel metal2 23632 24136 23632 24136 0 _088_
rlabel metal2 26040 18536 26040 18536 0 _089_
rlabel metal2 26376 22064 26376 22064 0 _090_
rlabel metal2 22120 23128 22120 23128 0 _091_
rlabel metal2 25704 21784 25704 21784 0 _092_
rlabel metal2 23016 20104 23016 20104 0 _093_
rlabel metal3 18256 17416 18256 17416 0 _094_
rlabel metal3 19768 17528 19768 17528 0 _095_
rlabel metal2 17528 19824 17528 19824 0 _096_
rlabel metal2 15624 19936 15624 19936 0 _097_
rlabel metal2 16912 27720 16912 27720 0 _098_
rlabel metal2 17640 27356 17640 27356 0 _099_
rlabel metal2 14000 26936 14000 26936 0 _100_
rlabel metal3 16632 27832 16632 27832 0 _101_
rlabel metal3 24640 27832 24640 27832 0 _102_
rlabel metal3 17696 23016 17696 23016 0 _103_
rlabel metal2 22456 22848 22456 22848 0 _104_
rlabel metal2 19432 21728 19432 21728 0 clk
rlabel metal3 20720 21448 20720 21448 0 clknet_0_clk
rlabel metal3 23912 14504 23912 14504 0 clknet_1_0__leaf_clk
rlabel metal2 20216 27384 20216 27384 0 clknet_1_1__leaf_clk
rlabel metal2 16856 23968 16856 23968 0 dut58.count\[0\]
rlabel metal2 20552 27160 20552 27160 0 dut58.count\[1\]
rlabel metal2 22344 24752 22344 24752 0 dut58.count\[2\]
rlabel metal2 23464 23128 23464 23128 0 dut58.count\[3\]
rlabel metal2 10024 19656 10024 19656 0 net1
rlabel metal2 12040 18760 12040 18760 0 net10
rlabel metal3 30716 20552 30716 20552 0 net11
rlabel metal2 29176 20832 29176 20832 0 net12
rlabel metal3 23800 27720 23800 27720 0 net13
rlabel metal2 14728 27888 14728 27888 0 net14
rlabel metal2 11368 27384 11368 27384 0 net15
rlabel metal2 17416 6356 17416 6356 0 net16
rlabel metal3 7616 23016 7616 23016 0 net17
rlabel metal2 25928 27608 25928 27608 0 net18
rlabel metal2 20776 16408 20776 16408 0 net19
rlabel metal3 31920 19096 31920 19096 0 net2
rlabel metal2 13496 16912 13496 16912 0 net20
rlabel metal2 21448 5964 21448 5964 0 net21
rlabel metal2 28728 25032 28728 25032 0 net22
rlabel metal2 28392 26600 28392 26600 0 net23
rlabel metal2 17528 29540 17528 29540 0 net24
rlabel metal2 40264 21280 40264 21280 0 net25
rlabel metal2 18200 1246 18200 1246 0 net26
rlabel metal2 25144 14168 25144 14168 0 net3
rlabel metal3 7504 21448 7504 21448 0 net4
rlabel metal2 27944 16856 27944 16856 0 net5
rlabel metal2 27944 6356 27944 6356 0 net6
rlabel metal2 28280 17304 28280 17304 0 net7
rlabel metal2 22120 13552 22120 13552 0 net8
rlabel metal2 17640 5964 17640 5964 0 net9
rlabel metal3 1358 19544 1358 19544 0 segm[10]
rlabel metal2 40040 19096 40040 19096 0 segm[11]
rlabel metal2 24920 2198 24920 2198 0 segm[12]
rlabel metal3 1358 21560 1358 21560 0 segm[13]
rlabel metal2 40040 17640 40040 17640 0 segm[1]
rlabel metal2 25592 2422 25592 2422 0 segm[2]
rlabel metal3 40642 18200 40642 18200 0 segm[4]
rlabel metal2 20888 2422 20888 2422 0 segm[5]
rlabel metal2 17528 2198 17528 2198 0 segm[6]
rlabel metal3 1358 18872 1358 18872 0 segm[7]
rlabel metal2 40040 20552 40040 20552 0 segm[8]
rlabel metal2 40040 19656 40040 19656 0 segm[9]
rlabel metal2 22904 39746 22904 39746 0 sel[0]
rlabel metal3 1358 27608 1358 27608 0 sel[10]
rlabel metal3 1358 26936 1358 26936 0 sel[11]
rlabel metal2 16856 2422 16856 2422 0 sel[1]
rlabel metal3 1358 23576 1358 23576 0 sel[2]
rlabel metal2 25592 39914 25592 39914 0 sel[3]
rlabel metal2 20216 2982 20216 2982 0 sel[4]
rlabel metal3 1358 16856 1358 16856 0 sel[5]
rlabel metal2 21560 2198 21560 2198 0 sel[6]
rlabel metal2 40040 25256 40040 25256 0 sel[7]
rlabel metal2 40040 27048 40040 27048 0 sel[8]
rlabel metal2 18200 39746 18200 39746 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
