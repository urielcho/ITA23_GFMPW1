magic
tech gf180mcuD
magscale 1 5
timestamp 1699643231
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9417 19055 9423 19081
rect 9449 19055 9455 19081
rect 9865 18999 9871 19025
rect 9897 18999 9903 19025
rect 10817 18999 10823 19025
rect 10849 18999 10855 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 14239 18969 14265 18975
rect 14239 18937 14265 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10711 18745 10737 18751
rect 10711 18713 10737 18719
rect 13399 18745 13425 18751
rect 13399 18713 13425 18719
rect 10201 18607 10207 18633
rect 10233 18607 10239 18633
rect 12889 18607 12895 18633
rect 12921 18607 12927 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 9815 14209 9841 14215
rect 9815 14177 9841 14183
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 9479 14041 9505 14047
rect 9479 14009 9505 14015
rect 8975 13985 9001 13991
rect 8975 13953 9001 13959
rect 8863 13929 8889 13935
rect 8863 13897 8889 13903
rect 9031 13929 9057 13935
rect 9031 13897 9057 13903
rect 9367 13929 9393 13935
rect 9367 13897 9393 13903
rect 9535 13929 9561 13935
rect 9865 13903 9871 13929
rect 9897 13903 9903 13929
rect 9535 13897 9561 13903
rect 11551 13873 11577 13879
rect 10257 13847 10263 13873
rect 10289 13847 10295 13873
rect 11321 13847 11327 13873
rect 11353 13847 11359 13873
rect 11551 13841 11577 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 9871 13649 9897 13655
rect 9871 13617 9897 13623
rect 10319 13649 10345 13655
rect 10319 13617 10345 13623
rect 967 13593 993 13599
rect 8577 13567 8583 13593
rect 8609 13567 8615 13593
rect 9641 13567 9647 13593
rect 9673 13567 9679 13593
rect 967 13561 993 13567
rect 2137 13511 2143 13537
rect 2169 13511 2175 13537
rect 8185 13511 8191 13537
rect 8217 13511 8223 13537
rect 7575 13481 7601 13487
rect 7575 13449 7601 13455
rect 7631 13481 7657 13487
rect 7631 13449 7657 13455
rect 9815 13481 9841 13487
rect 9815 13449 9841 13455
rect 9871 13481 9897 13487
rect 9871 13449 9897 13455
rect 10375 13481 10401 13487
rect 10375 13449 10401 13455
rect 10711 13481 10737 13487
rect 10711 13449 10737 13455
rect 10823 13481 10849 13487
rect 10823 13449 10849 13455
rect 10879 13481 10905 13487
rect 10879 13449 10905 13455
rect 7127 13425 7153 13431
rect 7127 13393 7153 13399
rect 7239 13425 7265 13431
rect 7239 13393 7265 13399
rect 7295 13425 7321 13431
rect 7295 13393 7321 13399
rect 7351 13425 7377 13431
rect 7351 13393 7377 13399
rect 7463 13425 7489 13431
rect 7463 13393 7489 13399
rect 10319 13425 10345 13431
rect 10319 13393 10345 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7631 13257 7657 13263
rect 7631 13225 7657 13231
rect 7743 13201 7769 13207
rect 7743 13169 7769 13175
rect 7799 13201 7825 13207
rect 7799 13169 7825 13175
rect 12671 13201 12697 13207
rect 12671 13169 12697 13175
rect 8023 13145 8049 13151
rect 11775 13145 11801 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 7513 13119 7519 13145
rect 7545 13119 7551 13145
rect 8689 13119 8695 13145
rect 8721 13119 8727 13145
rect 11657 13119 11663 13145
rect 11689 13119 11695 13145
rect 8023 13113 8049 13119
rect 11775 13113 11801 13119
rect 11887 13145 11913 13151
rect 12615 13145 12641 13151
rect 11993 13119 11999 13145
rect 12025 13119 12031 13145
rect 11887 13113 11913 13119
rect 12615 13113 12641 13119
rect 10375 13089 10401 13095
rect 6057 13063 6063 13089
rect 6089 13063 6095 13089
rect 7121 13063 7127 13089
rect 7153 13063 7159 13089
rect 9081 13063 9087 13089
rect 9113 13063 9119 13089
rect 10145 13063 10151 13089
rect 10177 13063 10183 13089
rect 10375 13057 10401 13063
rect 11831 13089 11857 13095
rect 11831 13057 11857 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 9367 12809 9393 12815
rect 11825 12783 11831 12809
rect 11857 12783 11863 12809
rect 12889 12783 12895 12809
rect 12921 12783 12927 12809
rect 9367 12777 9393 12783
rect 7575 12753 7601 12759
rect 7575 12721 7601 12727
rect 7687 12753 7713 12759
rect 7687 12721 7713 12727
rect 9647 12753 9673 12759
rect 9809 12727 9815 12753
rect 9841 12727 9847 12753
rect 11489 12727 11495 12753
rect 11521 12727 11527 12753
rect 13281 12727 13287 12753
rect 13313 12727 13319 12753
rect 9647 12721 9673 12727
rect 7295 12697 7321 12703
rect 7295 12665 7321 12671
rect 7407 12697 7433 12703
rect 7407 12665 7433 12671
rect 7463 12697 7489 12703
rect 13455 12697 13481 12703
rect 9921 12671 9927 12697
rect 9953 12671 9959 12697
rect 7463 12665 7489 12671
rect 13455 12665 13481 12671
rect 9311 12641 9337 12647
rect 9311 12609 9337 12615
rect 9423 12641 9449 12647
rect 9423 12609 9449 12615
rect 11271 12641 11297 12647
rect 11271 12609 11297 12615
rect 13119 12641 13145 12647
rect 13119 12609 13145 12615
rect 13399 12641 13425 12647
rect 13399 12609 13425 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 9249 12447 9255 12473
rect 9281 12447 9287 12473
rect 7233 12391 7239 12417
rect 7265 12391 7271 12417
rect 13393 12391 13399 12417
rect 13425 12391 13431 12417
rect 9423 12361 9449 12367
rect 7625 12335 7631 12361
rect 7657 12335 7663 12361
rect 9809 12335 9815 12361
rect 9841 12335 9847 12361
rect 13001 12335 13007 12361
rect 13033 12335 13039 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 9423 12329 9449 12335
rect 7855 12305 7881 12311
rect 12671 12305 12697 12311
rect 6169 12279 6175 12305
rect 6201 12279 6207 12305
rect 12105 12279 12111 12305
rect 12137 12279 12143 12305
rect 14457 12279 14463 12305
rect 14489 12279 14495 12305
rect 7855 12273 7881 12279
rect 12671 12273 12697 12279
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 967 12025 993 12031
rect 967 11993 993 11999
rect 8919 12025 8945 12031
rect 13959 12025 13985 12031
rect 12105 11999 12111 12025
rect 12137 11999 12143 12025
rect 13729 11999 13735 12025
rect 13761 11999 13767 12025
rect 8919 11993 8945 11999
rect 13959 11993 13985 11999
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 6903 11969 6929 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 6903 11937 6929 11943
rect 8415 11969 8441 11975
rect 10033 11943 10039 11969
rect 10065 11943 10071 11969
rect 10705 11943 10711 11969
rect 10737 11943 10743 11969
rect 12273 11943 12279 11969
rect 12305 11943 12311 11969
rect 14065 11943 14071 11969
rect 14097 11943 14103 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 8415 11937 8441 11943
rect 8583 11913 8609 11919
rect 8583 11881 8609 11887
rect 8695 11913 8721 11919
rect 8695 11881 8721 11887
rect 9871 11913 9897 11919
rect 9871 11881 9897 11887
rect 9927 11913 9953 11919
rect 13903 11913 13929 11919
rect 11041 11887 11047 11913
rect 11073 11887 11079 11913
rect 12665 11887 12671 11913
rect 12697 11887 12703 11913
rect 9927 11881 9953 11887
rect 13903 11881 13929 11887
rect 8471 11857 8497 11863
rect 8471 11825 8497 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 11047 11689 11073 11695
rect 11047 11657 11073 11663
rect 12783 11689 12809 11695
rect 12783 11657 12809 11663
rect 8695 11633 8721 11639
rect 8017 11607 8023 11633
rect 8049 11607 8055 11633
rect 8695 11601 8721 11607
rect 12055 11633 12081 11639
rect 12055 11601 12081 11607
rect 12279 11633 12305 11639
rect 12279 11601 12305 11607
rect 12839 11633 12865 11639
rect 12839 11601 12865 11607
rect 9535 11577 9561 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 6785 11551 6791 11577
rect 6817 11551 6823 11577
rect 8409 11551 8415 11577
rect 8441 11551 8447 11577
rect 8801 11551 8807 11577
rect 8833 11551 8839 11577
rect 9305 11551 9311 11577
rect 9337 11551 9343 11577
rect 9535 11545 9561 11551
rect 10207 11577 10233 11583
rect 10207 11545 10233 11551
rect 10319 11577 10345 11583
rect 10319 11545 10345 11551
rect 10543 11577 10569 11583
rect 10543 11545 10569 11551
rect 10599 11577 10625 11583
rect 10991 11577 11017 11583
rect 10761 11551 10767 11577
rect 10793 11551 10799 11577
rect 10599 11545 10625 11551
rect 10991 11545 11017 11551
rect 11103 11577 11129 11583
rect 11831 11577 11857 11583
rect 12895 11577 12921 11583
rect 11601 11551 11607 11577
rect 11633 11551 11639 11577
rect 12161 11551 12167 11577
rect 12193 11551 12199 11577
rect 12609 11551 12615 11577
rect 12641 11551 12647 11577
rect 11103 11545 11129 11551
rect 11831 11545 11857 11551
rect 12895 11545 12921 11551
rect 10039 11521 10065 11527
rect 5329 11495 5335 11521
rect 5361 11495 5367 11521
rect 6393 11495 6399 11521
rect 6425 11495 6431 11521
rect 6953 11495 6959 11521
rect 6985 11495 6991 11521
rect 10039 11489 10065 11495
rect 10263 11521 10289 11527
rect 10263 11489 10289 11495
rect 11495 11521 11521 11527
rect 12329 11495 12335 11521
rect 12361 11495 12367 11521
rect 11495 11489 11521 11495
rect 967 11465 993 11471
rect 9927 11465 9953 11471
rect 8857 11439 8863 11465
rect 8889 11439 8895 11465
rect 9753 11439 9759 11465
rect 9785 11439 9791 11465
rect 967 11433 993 11439
rect 9927 11433 9953 11439
rect 10879 11465 10905 11471
rect 10879 11433 10905 11439
rect 11439 11465 11465 11471
rect 11439 11433 11465 11439
rect 11887 11465 11913 11471
rect 11887 11433 11913 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 7687 11297 7713 11303
rect 7687 11265 7713 11271
rect 7911 11297 7937 11303
rect 7911 11265 7937 11271
rect 7967 11297 7993 11303
rect 7967 11265 7993 11271
rect 967 11241 993 11247
rect 967 11209 993 11215
rect 8751 11241 8777 11247
rect 8751 11209 8777 11215
rect 10151 11241 10177 11247
rect 11657 11215 11663 11241
rect 11689 11215 11695 11241
rect 10151 11209 10177 11215
rect 7799 11185 7825 11191
rect 8807 11185 8833 11191
rect 10263 11185 10289 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 8577 11159 8583 11185
rect 8609 11159 8615 11185
rect 9193 11159 9199 11185
rect 9225 11159 9231 11185
rect 10649 11159 10655 11185
rect 10681 11159 10687 11185
rect 11153 11159 11159 11185
rect 11185 11159 11191 11185
rect 11601 11159 11607 11185
rect 11633 11159 11639 11185
rect 7799 11153 7825 11159
rect 8807 11153 8833 11159
rect 10263 11153 10289 11159
rect 6735 11129 6761 11135
rect 6735 11097 6761 11103
rect 6903 11129 6929 11135
rect 6903 11097 6929 11103
rect 7631 11129 7657 11135
rect 7631 11097 7657 11103
rect 10095 11129 10121 11135
rect 10095 11097 10121 11103
rect 10375 11129 10401 11135
rect 11321 11103 11327 11129
rect 11353 11103 11359 11129
rect 11545 11103 11551 11129
rect 11577 11103 11583 11129
rect 10375 11097 10401 11103
rect 8695 11073 8721 11079
rect 8695 11041 8721 11047
rect 8863 11073 8889 11079
rect 12111 11073 12137 11079
rect 9081 11047 9087 11073
rect 9113 11047 9119 11073
rect 8863 11041 8889 11047
rect 12111 11041 12137 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 6959 10905 6985 10911
rect 6959 10873 6985 10879
rect 7799 10905 7825 10911
rect 7799 10873 7825 10879
rect 8919 10905 8945 10911
rect 9081 10879 9087 10905
rect 9113 10879 9119 10905
rect 12105 10879 12111 10905
rect 12137 10879 12143 10905
rect 8919 10873 8945 10879
rect 7239 10849 7265 10855
rect 7239 10817 7265 10823
rect 7351 10849 7377 10855
rect 7351 10817 7377 10823
rect 7407 10849 7433 10855
rect 7407 10817 7433 10823
rect 7631 10849 7657 10855
rect 7631 10817 7657 10823
rect 8807 10849 8833 10855
rect 8807 10817 8833 10823
rect 9591 10849 9617 10855
rect 11943 10849 11969 10855
rect 10369 10823 10375 10849
rect 10401 10823 10407 10849
rect 10929 10823 10935 10849
rect 10961 10823 10967 10849
rect 9591 10817 9617 10823
rect 11943 10817 11969 10823
rect 13231 10849 13257 10855
rect 13231 10817 13257 10823
rect 6847 10793 6873 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 6673 10767 6679 10793
rect 6705 10767 6711 10793
rect 6847 10761 6873 10767
rect 7183 10793 7209 10799
rect 7183 10761 7209 10767
rect 7743 10793 7769 10799
rect 7743 10761 7769 10767
rect 7855 10793 7881 10799
rect 8751 10793 8777 10799
rect 9703 10793 9729 10799
rect 12727 10793 12753 10799
rect 13063 10793 13089 10799
rect 7961 10767 7967 10793
rect 7993 10767 7999 10793
rect 9193 10767 9199 10793
rect 9225 10767 9231 10793
rect 11265 10767 11271 10793
rect 11297 10767 11303 10793
rect 11713 10767 11719 10793
rect 11745 10767 11751 10793
rect 12217 10767 12223 10793
rect 12249 10767 12255 10793
rect 12889 10767 12895 10793
rect 12921 10767 12927 10793
rect 7855 10761 7881 10767
rect 8751 10761 8777 10767
rect 9703 10761 9729 10767
rect 12727 10761 12753 10767
rect 13063 10761 13089 10767
rect 967 10737 993 10743
rect 6903 10737 6929 10743
rect 12615 10737 12641 10743
rect 5217 10711 5223 10737
rect 5249 10711 5255 10737
rect 6281 10711 6287 10737
rect 6313 10711 6319 10737
rect 11489 10711 11495 10737
rect 11521 10711 11527 10737
rect 967 10705 993 10711
rect 6903 10705 6929 10711
rect 12615 10705 12641 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 11153 10487 11159 10513
rect 11185 10487 11191 10513
rect 7127 10457 7153 10463
rect 11215 10457 11241 10463
rect 8633 10431 8639 10457
rect 8665 10431 8671 10457
rect 11881 10431 11887 10457
rect 11913 10431 11919 10457
rect 13225 10431 13231 10457
rect 13257 10431 13263 10457
rect 14289 10431 14295 10457
rect 14321 10431 14327 10457
rect 7127 10425 7153 10431
rect 11215 10425 11241 10431
rect 6903 10401 6929 10407
rect 9087 10401 9113 10407
rect 8801 10375 8807 10401
rect 8833 10375 8839 10401
rect 6903 10369 6929 10375
rect 9087 10369 9113 10375
rect 9871 10401 9897 10407
rect 11607 10401 11633 10407
rect 12279 10401 12305 10407
rect 10593 10375 10599 10401
rect 10625 10375 10631 10401
rect 10985 10375 10991 10401
rect 11017 10375 11023 10401
rect 11769 10375 11775 10401
rect 11801 10375 11807 10401
rect 9871 10369 9897 10375
rect 11607 10369 11633 10375
rect 12279 10369 12305 10375
rect 12559 10401 12585 10407
rect 12889 10375 12895 10401
rect 12921 10375 12927 10401
rect 12559 10369 12585 10375
rect 9031 10345 9057 10351
rect 6729 10319 6735 10345
rect 6761 10319 6767 10345
rect 10033 10319 10039 10345
rect 10065 10319 10071 10345
rect 9031 10313 9057 10319
rect 9479 10289 9505 10295
rect 9479 10257 9505 10263
rect 11439 10289 11465 10295
rect 11439 10257 11465 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 12951 10121 12977 10127
rect 12951 10089 12977 10095
rect 8023 10065 8049 10071
rect 6337 10039 6343 10065
rect 6369 10039 6375 10065
rect 8023 10033 8049 10039
rect 8359 10065 8385 10071
rect 8359 10033 8385 10039
rect 8863 10065 8889 10071
rect 8863 10033 8889 10039
rect 9199 10065 9225 10071
rect 12671 10065 12697 10071
rect 10929 10039 10935 10065
rect 10961 10039 10967 10065
rect 9199 10033 9225 10039
rect 12671 10033 12697 10039
rect 8247 10009 8273 10015
rect 6001 9983 6007 10009
rect 6033 9983 6039 10009
rect 8247 9977 8273 9983
rect 8415 10009 8441 10015
rect 8415 9977 8441 9983
rect 8695 10009 8721 10015
rect 9641 9983 9647 10009
rect 9673 9983 9679 10009
rect 13113 9983 13119 10009
rect 13145 9983 13151 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 8695 9977 8721 9983
rect 7687 9953 7713 9959
rect 7401 9927 7407 9953
rect 7433 9927 7439 9953
rect 7687 9921 7713 9927
rect 12615 9953 12641 9959
rect 13505 9927 13511 9953
rect 13537 9927 13543 9953
rect 14569 9927 14575 9953
rect 14601 9927 14607 9953
rect 12615 9921 12641 9927
rect 7967 9897 7993 9903
rect 7967 9865 7993 9871
rect 8135 9897 8161 9903
rect 8135 9865 8161 9871
rect 9311 9897 9337 9903
rect 9311 9865 9337 9871
rect 9479 9897 9505 9903
rect 9479 9865 9505 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8415 9729 8441 9735
rect 10207 9729 10233 9735
rect 8745 9703 8751 9729
rect 8777 9703 8783 9729
rect 8415 9697 8441 9703
rect 10207 9697 10233 9703
rect 11999 9729 12025 9735
rect 13505 9703 13511 9729
rect 13537 9703 13543 9729
rect 11999 9697 12025 9703
rect 10263 9673 10289 9679
rect 9417 9647 9423 9673
rect 9449 9647 9455 9673
rect 10263 9641 10289 9647
rect 10711 9673 10737 9679
rect 10711 9641 10737 9647
rect 13847 9673 13873 9679
rect 13847 9641 13873 9647
rect 6903 9617 6929 9623
rect 6903 9585 6929 9591
rect 8919 9617 8945 9623
rect 8919 9585 8945 9591
rect 9031 9617 9057 9623
rect 10599 9617 10625 9623
rect 9249 9591 9255 9617
rect 9281 9591 9287 9617
rect 9031 9585 9057 9591
rect 10599 9585 10625 9591
rect 10879 9617 10905 9623
rect 10879 9585 10905 9591
rect 11327 9617 11353 9623
rect 11327 9585 11353 9591
rect 11551 9617 11577 9623
rect 12223 9617 12249 9623
rect 11769 9591 11775 9617
rect 11801 9591 11807 9617
rect 11551 9585 11577 9591
rect 12223 9585 12249 9591
rect 12503 9617 12529 9623
rect 12503 9585 12529 9591
rect 13231 9617 13257 9623
rect 13617 9591 13623 9617
rect 13649 9591 13655 9617
rect 13953 9591 13959 9617
rect 13985 9591 13991 9617
rect 13231 9585 13257 9591
rect 6735 9561 6761 9567
rect 6735 9529 6761 9535
rect 8471 9561 8497 9567
rect 8471 9529 8497 9535
rect 8583 9561 8609 9567
rect 8583 9529 8609 9535
rect 10319 9561 10345 9567
rect 10319 9529 10345 9535
rect 10823 9561 10849 9567
rect 13791 9561 13817 9567
rect 12049 9535 12055 9561
rect 12081 9535 12087 9561
rect 13337 9535 13343 9561
rect 13369 9535 13375 9561
rect 10823 9529 10849 9535
rect 13791 9529 13817 9535
rect 9647 9505 9673 9511
rect 11495 9505 11521 9511
rect 9809 9479 9815 9505
rect 9841 9479 9847 9505
rect 9647 9473 9673 9479
rect 11495 9473 11521 9479
rect 12951 9505 12977 9511
rect 13449 9479 13455 9505
rect 13481 9479 13487 9505
rect 12951 9473 12977 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 9311 9337 9337 9343
rect 9025 9311 9031 9337
rect 9057 9311 9063 9337
rect 9311 9305 9337 9311
rect 10151 9337 10177 9343
rect 10151 9305 10177 9311
rect 10263 9337 10289 9343
rect 10263 9305 10289 9311
rect 11327 9337 11353 9343
rect 12777 9311 12783 9337
rect 12809 9311 12815 9337
rect 11327 9305 11353 9311
rect 10095 9281 10121 9287
rect 9753 9255 9759 9281
rect 9785 9255 9791 9281
rect 11601 9255 11607 9281
rect 11633 9255 11639 9281
rect 10095 9249 10121 9255
rect 7015 9225 7041 9231
rect 7015 9193 7041 9199
rect 7183 9225 7209 9231
rect 7183 9193 7209 9199
rect 7351 9225 7377 9231
rect 9143 9225 9169 9231
rect 8913 9199 8919 9225
rect 8945 9199 8951 9225
rect 7351 9193 7377 9199
rect 9143 9193 9169 9199
rect 9311 9225 9337 9231
rect 9311 9193 9337 9199
rect 9479 9225 9505 9231
rect 11103 9225 11129 9231
rect 9865 9199 9871 9225
rect 9897 9199 9903 9225
rect 9479 9193 9505 9199
rect 11103 9193 11129 9199
rect 11439 9225 11465 9231
rect 11439 9193 11465 9199
rect 11775 9225 11801 9231
rect 11775 9193 11801 9199
rect 12615 9225 12641 9231
rect 12615 9193 12641 9199
rect 7127 9169 7153 9175
rect 10873 9143 10879 9169
rect 10905 9143 10911 9169
rect 11265 9143 11271 9169
rect 11297 9143 11303 9169
rect 7127 9137 7153 9143
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 11383 8945 11409 8951
rect 11383 8913 11409 8919
rect 967 8889 993 8895
rect 967 8857 993 8863
rect 8975 8889 9001 8895
rect 8975 8857 9001 8863
rect 9479 8889 9505 8895
rect 9479 8857 9505 8863
rect 10319 8889 10345 8895
rect 10319 8857 10345 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 8527 8833 8553 8839
rect 9815 8833 9841 8839
rect 12055 8833 12081 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 8801 8807 8807 8833
rect 8833 8807 8839 8833
rect 9361 8807 9367 8833
rect 9393 8807 9399 8833
rect 10649 8807 10655 8833
rect 10681 8807 10687 8833
rect 11153 8807 11159 8833
rect 11185 8807 11191 8833
rect 11881 8807 11887 8833
rect 11913 8807 11919 8833
rect 12385 8807 12391 8833
rect 12417 8807 12423 8833
rect 13225 8807 13231 8833
rect 13257 8807 13263 8833
rect 18937 8807 18943 8833
rect 18969 8807 18975 8833
rect 8527 8801 8553 8807
rect 9815 8801 9841 8807
rect 12055 8801 12081 8807
rect 9535 8777 9561 8783
rect 9535 8745 9561 8751
rect 10263 8777 10289 8783
rect 11439 8777 11465 8783
rect 10705 8751 10711 8777
rect 10737 8751 10743 8777
rect 10263 8745 10289 8751
rect 11439 8745 11465 8751
rect 11607 8777 11633 8783
rect 11607 8745 11633 8751
rect 13399 8777 13425 8783
rect 13399 8745 13425 8751
rect 8751 8721 8777 8727
rect 8353 8695 8359 8721
rect 8385 8695 8391 8721
rect 8751 8689 8777 8695
rect 9871 8721 9897 8727
rect 9871 8689 9897 8695
rect 9983 8721 10009 8727
rect 9983 8689 10009 8695
rect 10151 8721 10177 8727
rect 10151 8689 10177 8695
rect 10375 8721 10401 8727
rect 13343 8721 13369 8727
rect 11153 8695 11159 8721
rect 11185 8695 11191 8721
rect 12273 8695 12279 8721
rect 12305 8695 12311 8721
rect 10375 8689 10401 8695
rect 13343 8689 13369 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7295 8553 7321 8559
rect 7295 8521 7321 8527
rect 7575 8553 7601 8559
rect 7575 8521 7601 8527
rect 8807 8553 8833 8559
rect 8807 8521 8833 8527
rect 8863 8497 8889 8503
rect 13337 8471 13343 8497
rect 13369 8471 13375 8497
rect 8863 8465 8889 8471
rect 7239 8441 7265 8447
rect 12783 8441 12809 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7009 8415 7015 8441
rect 7041 8415 7047 8441
rect 9697 8415 9703 8441
rect 9729 8415 9735 8441
rect 11377 8415 11383 8441
rect 11409 8415 11415 8441
rect 12945 8415 12951 8441
rect 12977 8415 12983 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 7239 8409 7265 8415
rect 12783 8409 12809 8415
rect 5609 8359 5615 8385
rect 5641 8359 5647 8385
rect 6673 8359 6679 8385
rect 6705 8359 6711 8385
rect 14401 8359 14407 8385
rect 14433 8359 14439 8385
rect 19945 8359 19951 8385
rect 19977 8359 19983 8385
rect 967 8329 993 8335
rect 967 8297 993 8303
rect 7295 8329 7321 8335
rect 7295 8297 7321 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 6455 8161 6481 8167
rect 6455 8129 6481 8135
rect 6959 8161 6985 8167
rect 6959 8129 6985 8135
rect 12055 8161 12081 8167
rect 12055 8129 12081 8135
rect 13175 8161 13201 8167
rect 13175 8129 13201 8135
rect 6399 8105 6425 8111
rect 13623 8105 13649 8111
rect 7905 8079 7911 8105
rect 7937 8079 7943 8105
rect 8969 8079 8975 8105
rect 9001 8079 9007 8105
rect 12721 8079 12727 8105
rect 12753 8079 12759 8105
rect 6399 8073 6425 8079
rect 13623 8073 13649 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 10263 8049 10289 8055
rect 7569 8023 7575 8049
rect 7601 8023 7607 8049
rect 10263 8017 10289 8023
rect 10655 8049 10681 8055
rect 10655 8017 10681 8023
rect 10767 8049 10793 8055
rect 12503 8049 12529 8055
rect 13063 8049 13089 8055
rect 11265 8023 11271 8049
rect 11297 8023 11303 8049
rect 12105 8023 12111 8049
rect 12137 8023 12143 8049
rect 12945 8023 12951 8049
rect 12977 8023 12983 8049
rect 10767 8017 10793 8023
rect 12503 8017 12529 8023
rect 13063 8017 13089 8023
rect 13343 8049 13369 8055
rect 13343 8017 13369 8023
rect 13567 8049 13593 8055
rect 13567 8017 13593 8023
rect 13679 8049 13705 8055
rect 13679 8017 13705 8023
rect 13847 8049 13873 8055
rect 13847 8017 13873 8023
rect 13903 8049 13929 8055
rect 14009 8023 14015 8049
rect 14041 8023 14047 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 13903 8017 13929 8023
rect 7015 7993 7041 7999
rect 7015 7961 7041 7967
rect 10319 7993 10345 7999
rect 10319 7961 10345 7967
rect 11159 7993 11185 7999
rect 11159 7961 11185 7967
rect 11495 7993 11521 7999
rect 11831 7993 11857 7999
rect 13231 7993 13257 7999
rect 11657 7967 11663 7993
rect 11689 7967 11695 7993
rect 11937 7967 11943 7993
rect 11969 7967 11975 7993
rect 11495 7961 11521 7967
rect 11831 7961 11857 7967
rect 13231 7961 13257 7967
rect 6959 7937 6985 7943
rect 6959 7905 6985 7911
rect 9199 7937 9225 7943
rect 9199 7905 9225 7911
rect 10431 7937 10457 7943
rect 10431 7905 10457 7911
rect 10711 7937 10737 7943
rect 10711 7905 10737 7911
rect 10879 7937 10905 7943
rect 10879 7905 10905 7911
rect 11887 7937 11913 7943
rect 11887 7905 11913 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 7575 7769 7601 7775
rect 7575 7737 7601 7743
rect 8919 7769 8945 7775
rect 8919 7737 8945 7743
rect 9927 7769 9953 7775
rect 9927 7737 9953 7743
rect 10039 7769 10065 7775
rect 10039 7737 10065 7743
rect 12895 7769 12921 7775
rect 12895 7737 12921 7743
rect 8863 7713 8889 7719
rect 6953 7687 6959 7713
rect 6985 7687 6991 7713
rect 8863 7681 8889 7687
rect 9031 7713 9057 7719
rect 9031 7681 9057 7687
rect 9815 7713 9841 7719
rect 13449 7687 13455 7713
rect 13481 7687 13487 7713
rect 14849 7687 14855 7713
rect 14881 7687 14887 7713
rect 9815 7681 9841 7687
rect 8751 7657 8777 7663
rect 7345 7631 7351 7657
rect 7377 7631 7383 7657
rect 8751 7625 8777 7631
rect 8807 7657 8833 7663
rect 8807 7625 8833 7631
rect 11607 7657 11633 7663
rect 11607 7625 11633 7631
rect 11775 7657 11801 7663
rect 11775 7625 11801 7631
rect 11887 7657 11913 7663
rect 13057 7631 13063 7657
rect 13089 7631 13095 7657
rect 14737 7631 14743 7657
rect 14769 7631 14775 7657
rect 18825 7631 18831 7657
rect 18857 7631 18863 7657
rect 11887 7625 11913 7631
rect 9983 7601 10009 7607
rect 5889 7575 5895 7601
rect 5921 7575 5927 7601
rect 9983 7569 10009 7575
rect 11719 7601 11745 7607
rect 20007 7601 20033 7607
rect 14513 7575 14519 7601
rect 14545 7575 14551 7601
rect 11719 7569 11745 7575
rect 20007 7569 20033 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9815 7377 9841 7383
rect 9815 7345 9841 7351
rect 9255 7321 9281 7327
rect 13287 7321 13313 7327
rect 9025 7295 9031 7321
rect 9057 7295 9063 7321
rect 11657 7295 11663 7321
rect 11689 7295 11695 7321
rect 12721 7295 12727 7321
rect 12753 7295 12759 7321
rect 9255 7289 9281 7295
rect 13287 7289 13313 7295
rect 7569 7239 7575 7265
rect 7601 7239 7607 7265
rect 11321 7239 11327 7265
rect 11353 7239 11359 7265
rect 14625 7239 14631 7265
rect 14657 7239 14663 7265
rect 7961 7183 7967 7209
rect 7993 7183 7999 7209
rect 9871 7181 9897 7187
rect 9815 7153 9841 7159
rect 9871 7149 9897 7155
rect 12895 7153 12921 7159
rect 9815 7121 9841 7127
rect 13057 7127 13063 7153
rect 13089 7127 13095 7153
rect 14737 7127 14743 7153
rect 14769 7127 14775 7153
rect 12895 7121 12921 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8359 6985 8385 6991
rect 8359 6953 8385 6959
rect 11775 6985 11801 6991
rect 11775 6953 11801 6959
rect 8415 6929 8441 6935
rect 10481 6903 10487 6929
rect 10513 6903 10519 6929
rect 8415 6897 8441 6903
rect 10145 6847 10151 6873
rect 10177 6847 10183 6873
rect 11545 6791 11551 6817
rect 11577 6791 11583 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 10767 6537 10793 6543
rect 9249 6511 9255 6537
rect 9281 6511 9287 6537
rect 10313 6511 10319 6537
rect 10345 6511 10351 6537
rect 10767 6505 10793 6511
rect 8913 6455 8919 6481
rect 8945 6455 8951 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 12889 2143 12895 2169
rect 12921 2143 12927 2169
rect 13399 2057 13425 2063
rect 13399 2025 13425 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 13063 1833 13089 1839
rect 13063 1801 13089 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10369 1751 10375 1777
rect 10401 1751 10407 1777
rect 12609 1751 12615 1777
rect 12641 1751 12647 1777
rect 10879 1665 10905 1671
rect 10879 1633 10905 1639
rect 12279 1665 12305 1671
rect 12279 1633 12305 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 9423 19055 9449 19081
rect 9871 18999 9897 19025
rect 10823 18999 10849 19025
rect 12279 18999 12305 19025
rect 14239 18943 14265 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10711 18719 10737 18745
rect 13399 18719 13425 18745
rect 10207 18607 10233 18633
rect 12895 18607 12921 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9815 14183 9841 14209
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 9479 14015 9505 14041
rect 8975 13959 9001 13985
rect 8863 13903 8889 13929
rect 9031 13903 9057 13929
rect 9367 13903 9393 13929
rect 9535 13903 9561 13929
rect 9871 13903 9897 13929
rect 10263 13847 10289 13873
rect 11327 13847 11353 13873
rect 11551 13847 11577 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9871 13623 9897 13649
rect 10319 13623 10345 13649
rect 967 13567 993 13593
rect 8583 13567 8609 13593
rect 9647 13567 9673 13593
rect 2143 13511 2169 13537
rect 8191 13511 8217 13537
rect 7575 13455 7601 13481
rect 7631 13455 7657 13481
rect 9815 13455 9841 13481
rect 9871 13455 9897 13481
rect 10375 13455 10401 13481
rect 10711 13455 10737 13481
rect 10823 13455 10849 13481
rect 10879 13455 10905 13481
rect 7127 13399 7153 13425
rect 7239 13399 7265 13425
rect 7295 13399 7321 13425
rect 7351 13399 7377 13425
rect 7463 13399 7489 13425
rect 10319 13399 10345 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7631 13231 7657 13257
rect 7743 13175 7769 13201
rect 7799 13175 7825 13201
rect 12671 13175 12697 13201
rect 2143 13119 2169 13145
rect 7519 13119 7545 13145
rect 8023 13119 8049 13145
rect 8695 13119 8721 13145
rect 11663 13119 11689 13145
rect 11775 13119 11801 13145
rect 11887 13119 11913 13145
rect 11999 13119 12025 13145
rect 12615 13119 12641 13145
rect 6063 13063 6089 13089
rect 7127 13063 7153 13089
rect 9087 13063 9113 13089
rect 10151 13063 10177 13089
rect 10375 13063 10401 13089
rect 11831 13063 11857 13089
rect 967 13007 993 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 9367 12783 9393 12809
rect 11831 12783 11857 12809
rect 12895 12783 12921 12809
rect 7575 12727 7601 12753
rect 7687 12727 7713 12753
rect 9647 12727 9673 12753
rect 9815 12727 9841 12753
rect 11495 12727 11521 12753
rect 13287 12727 13313 12753
rect 7295 12671 7321 12697
rect 7407 12671 7433 12697
rect 7463 12671 7489 12697
rect 9927 12671 9953 12697
rect 13455 12671 13481 12697
rect 9311 12615 9337 12641
rect 9423 12615 9449 12641
rect 11271 12615 11297 12641
rect 13119 12615 13145 12641
rect 13399 12615 13425 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 9255 12447 9281 12473
rect 7239 12391 7265 12417
rect 13399 12391 13425 12417
rect 7631 12335 7657 12361
rect 9423 12335 9449 12361
rect 9815 12335 9841 12361
rect 13007 12335 13033 12361
rect 18831 12335 18857 12361
rect 6175 12279 6201 12305
rect 7855 12279 7881 12305
rect 12111 12279 12137 12305
rect 12671 12279 12697 12305
rect 14463 12279 14489 12305
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 967 11999 993 12025
rect 8919 11999 8945 12025
rect 12111 11999 12137 12025
rect 13735 11999 13761 12025
rect 13959 11999 13985 12025
rect 20007 11999 20033 12025
rect 2143 11943 2169 11969
rect 6903 11943 6929 11969
rect 8415 11943 8441 11969
rect 10039 11943 10065 11969
rect 10711 11943 10737 11969
rect 12279 11943 12305 11969
rect 14071 11943 14097 11969
rect 18831 11943 18857 11969
rect 8583 11887 8609 11913
rect 8695 11887 8721 11913
rect 9871 11887 9897 11913
rect 9927 11887 9953 11913
rect 11047 11887 11073 11913
rect 12671 11887 12697 11913
rect 13903 11887 13929 11913
rect 8471 11831 8497 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 11047 11663 11073 11689
rect 12783 11663 12809 11689
rect 8023 11607 8049 11633
rect 8695 11607 8721 11633
rect 12055 11607 12081 11633
rect 12279 11607 12305 11633
rect 12839 11607 12865 11633
rect 2143 11551 2169 11577
rect 6791 11551 6817 11577
rect 8415 11551 8441 11577
rect 8807 11551 8833 11577
rect 9311 11551 9337 11577
rect 9535 11551 9561 11577
rect 10207 11551 10233 11577
rect 10319 11551 10345 11577
rect 10543 11551 10569 11577
rect 10599 11551 10625 11577
rect 10767 11551 10793 11577
rect 10991 11551 11017 11577
rect 11103 11551 11129 11577
rect 11607 11551 11633 11577
rect 11831 11551 11857 11577
rect 12167 11551 12193 11577
rect 12615 11551 12641 11577
rect 12895 11551 12921 11577
rect 5335 11495 5361 11521
rect 6399 11495 6425 11521
rect 6959 11495 6985 11521
rect 10039 11495 10065 11521
rect 10263 11495 10289 11521
rect 11495 11495 11521 11521
rect 12335 11495 12361 11521
rect 967 11439 993 11465
rect 8863 11439 8889 11465
rect 9759 11439 9785 11465
rect 9927 11439 9953 11465
rect 10879 11439 10905 11465
rect 11439 11439 11465 11465
rect 11887 11439 11913 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7687 11271 7713 11297
rect 7911 11271 7937 11297
rect 7967 11271 7993 11297
rect 967 11215 993 11241
rect 8751 11215 8777 11241
rect 10151 11215 10177 11241
rect 11663 11215 11689 11241
rect 2143 11159 2169 11185
rect 7799 11159 7825 11185
rect 8583 11159 8609 11185
rect 8807 11159 8833 11185
rect 9199 11159 9225 11185
rect 10263 11159 10289 11185
rect 10655 11159 10681 11185
rect 11159 11159 11185 11185
rect 11607 11159 11633 11185
rect 6735 11103 6761 11129
rect 6903 11103 6929 11129
rect 7631 11103 7657 11129
rect 10095 11103 10121 11129
rect 10375 11103 10401 11129
rect 11327 11103 11353 11129
rect 11551 11103 11577 11129
rect 8695 11047 8721 11073
rect 8863 11047 8889 11073
rect 9087 11047 9113 11073
rect 12111 11047 12137 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 6959 10879 6985 10905
rect 7799 10879 7825 10905
rect 8919 10879 8945 10905
rect 9087 10879 9113 10905
rect 12111 10879 12137 10905
rect 7239 10823 7265 10849
rect 7351 10823 7377 10849
rect 7407 10823 7433 10849
rect 7631 10823 7657 10849
rect 8807 10823 8833 10849
rect 9591 10823 9617 10849
rect 10375 10823 10401 10849
rect 10935 10823 10961 10849
rect 11943 10823 11969 10849
rect 13231 10823 13257 10849
rect 2143 10767 2169 10793
rect 6679 10767 6705 10793
rect 6847 10767 6873 10793
rect 7183 10767 7209 10793
rect 7743 10767 7769 10793
rect 7855 10767 7881 10793
rect 7967 10767 7993 10793
rect 8751 10767 8777 10793
rect 9199 10767 9225 10793
rect 9703 10767 9729 10793
rect 11271 10767 11297 10793
rect 11719 10767 11745 10793
rect 12223 10767 12249 10793
rect 12727 10767 12753 10793
rect 12895 10767 12921 10793
rect 13063 10767 13089 10793
rect 967 10711 993 10737
rect 5223 10711 5249 10737
rect 6287 10711 6313 10737
rect 6903 10711 6929 10737
rect 11495 10711 11521 10737
rect 12615 10711 12641 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 11159 10487 11185 10513
rect 7127 10431 7153 10457
rect 8639 10431 8665 10457
rect 11215 10431 11241 10457
rect 11887 10431 11913 10457
rect 13231 10431 13257 10457
rect 14295 10431 14321 10457
rect 6903 10375 6929 10401
rect 8807 10375 8833 10401
rect 9087 10375 9113 10401
rect 9871 10375 9897 10401
rect 10599 10375 10625 10401
rect 10991 10375 11017 10401
rect 11607 10375 11633 10401
rect 11775 10375 11801 10401
rect 12279 10375 12305 10401
rect 12559 10375 12585 10401
rect 12895 10375 12921 10401
rect 6735 10319 6761 10345
rect 9031 10319 9057 10345
rect 10039 10319 10065 10345
rect 9479 10263 9505 10289
rect 11439 10263 11465 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 12951 10095 12977 10121
rect 6343 10039 6369 10065
rect 8023 10039 8049 10065
rect 8359 10039 8385 10065
rect 8863 10039 8889 10065
rect 9199 10039 9225 10065
rect 10935 10039 10961 10065
rect 12671 10039 12697 10065
rect 6007 9983 6033 10009
rect 8247 9983 8273 10009
rect 8415 9983 8441 10009
rect 8695 9983 8721 10009
rect 9647 9983 9673 10009
rect 13119 9983 13145 10009
rect 18831 9983 18857 10009
rect 7407 9927 7433 9953
rect 7687 9927 7713 9953
rect 12615 9927 12641 9953
rect 13511 9927 13537 9953
rect 14575 9927 14601 9953
rect 7967 9871 7993 9897
rect 8135 9871 8161 9897
rect 9311 9871 9337 9897
rect 9479 9871 9505 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8415 9703 8441 9729
rect 8751 9703 8777 9729
rect 10207 9703 10233 9729
rect 11999 9703 12025 9729
rect 13511 9703 13537 9729
rect 9423 9647 9449 9673
rect 10263 9647 10289 9673
rect 10711 9647 10737 9673
rect 13847 9647 13873 9673
rect 6903 9591 6929 9617
rect 8919 9591 8945 9617
rect 9031 9591 9057 9617
rect 9255 9591 9281 9617
rect 10599 9591 10625 9617
rect 10879 9591 10905 9617
rect 11327 9591 11353 9617
rect 11551 9591 11577 9617
rect 11775 9591 11801 9617
rect 12223 9591 12249 9617
rect 12503 9591 12529 9617
rect 13231 9591 13257 9617
rect 13623 9591 13649 9617
rect 13959 9591 13985 9617
rect 6735 9535 6761 9561
rect 8471 9535 8497 9561
rect 8583 9535 8609 9561
rect 10319 9535 10345 9561
rect 10823 9535 10849 9561
rect 12055 9535 12081 9561
rect 13343 9535 13369 9561
rect 13791 9535 13817 9561
rect 9647 9479 9673 9505
rect 9815 9479 9841 9505
rect 11495 9479 11521 9505
rect 12951 9479 12977 9505
rect 13455 9479 13481 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 9031 9311 9057 9337
rect 9311 9311 9337 9337
rect 10151 9311 10177 9337
rect 10263 9311 10289 9337
rect 11327 9311 11353 9337
rect 12783 9311 12809 9337
rect 9759 9255 9785 9281
rect 10095 9255 10121 9281
rect 11607 9255 11633 9281
rect 7015 9199 7041 9225
rect 7183 9199 7209 9225
rect 7351 9199 7377 9225
rect 8919 9199 8945 9225
rect 9143 9199 9169 9225
rect 9311 9199 9337 9225
rect 9479 9199 9505 9225
rect 9871 9199 9897 9225
rect 11103 9199 11129 9225
rect 11439 9199 11465 9225
rect 11775 9199 11801 9225
rect 12615 9199 12641 9225
rect 7127 9143 7153 9169
rect 10879 9143 10905 9169
rect 11271 9143 11297 9169
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 11383 8919 11409 8945
rect 967 8863 993 8889
rect 8975 8863 9001 8889
rect 9479 8863 9505 8889
rect 10319 8863 10345 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 8527 8807 8553 8833
rect 8807 8807 8833 8833
rect 9367 8807 9393 8833
rect 9815 8807 9841 8833
rect 10655 8807 10681 8833
rect 11159 8807 11185 8833
rect 11887 8807 11913 8833
rect 12055 8807 12081 8833
rect 12391 8807 12417 8833
rect 13231 8807 13257 8833
rect 18943 8807 18969 8833
rect 9535 8751 9561 8777
rect 10263 8751 10289 8777
rect 10711 8751 10737 8777
rect 11439 8751 11465 8777
rect 11607 8751 11633 8777
rect 13399 8751 13425 8777
rect 8359 8695 8385 8721
rect 8751 8695 8777 8721
rect 9871 8695 9897 8721
rect 9983 8695 10009 8721
rect 10151 8695 10177 8721
rect 10375 8695 10401 8721
rect 11159 8695 11185 8721
rect 12279 8695 12305 8721
rect 13343 8695 13369 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7295 8527 7321 8553
rect 7575 8527 7601 8553
rect 8807 8527 8833 8553
rect 8863 8471 8889 8497
rect 13343 8471 13369 8497
rect 2143 8415 2169 8441
rect 7015 8415 7041 8441
rect 7239 8415 7265 8441
rect 9703 8415 9729 8441
rect 11383 8415 11409 8441
rect 12783 8415 12809 8441
rect 12951 8415 12977 8441
rect 18831 8415 18857 8441
rect 5615 8359 5641 8385
rect 6679 8359 6705 8385
rect 14407 8359 14433 8385
rect 19951 8359 19977 8385
rect 967 8303 993 8329
rect 7295 8303 7321 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 6455 8135 6481 8161
rect 6959 8135 6985 8161
rect 12055 8135 12081 8161
rect 13175 8135 13201 8161
rect 6399 8079 6425 8105
rect 7911 8079 7937 8105
rect 8975 8079 9001 8105
rect 12727 8079 12753 8105
rect 13623 8079 13649 8105
rect 20007 8079 20033 8105
rect 7575 8023 7601 8049
rect 10263 8023 10289 8049
rect 10655 8023 10681 8049
rect 10767 8023 10793 8049
rect 11271 8023 11297 8049
rect 12111 8023 12137 8049
rect 12503 8023 12529 8049
rect 12951 8023 12977 8049
rect 13063 8023 13089 8049
rect 13343 8023 13369 8049
rect 13567 8023 13593 8049
rect 13679 8023 13705 8049
rect 13847 8023 13873 8049
rect 13903 8023 13929 8049
rect 14015 8023 14041 8049
rect 18831 8023 18857 8049
rect 7015 7967 7041 7993
rect 10319 7967 10345 7993
rect 11159 7967 11185 7993
rect 11495 7967 11521 7993
rect 11663 7967 11689 7993
rect 11831 7967 11857 7993
rect 11943 7967 11969 7993
rect 13231 7967 13257 7993
rect 6959 7911 6985 7937
rect 9199 7911 9225 7937
rect 10431 7911 10457 7937
rect 10711 7911 10737 7937
rect 10879 7911 10905 7937
rect 11887 7911 11913 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 7575 7743 7601 7769
rect 8919 7743 8945 7769
rect 9927 7743 9953 7769
rect 10039 7743 10065 7769
rect 12895 7743 12921 7769
rect 6959 7687 6985 7713
rect 8863 7687 8889 7713
rect 9031 7687 9057 7713
rect 9815 7687 9841 7713
rect 13455 7687 13481 7713
rect 14855 7687 14881 7713
rect 7351 7631 7377 7657
rect 8751 7631 8777 7657
rect 8807 7631 8833 7657
rect 11607 7631 11633 7657
rect 11775 7631 11801 7657
rect 11887 7631 11913 7657
rect 13063 7631 13089 7657
rect 14743 7631 14769 7657
rect 18831 7631 18857 7657
rect 5895 7575 5921 7601
rect 9983 7575 10009 7601
rect 11719 7575 11745 7601
rect 14519 7575 14545 7601
rect 20007 7575 20033 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9815 7351 9841 7377
rect 9031 7295 9057 7321
rect 9255 7295 9281 7321
rect 11663 7295 11689 7321
rect 12727 7295 12753 7321
rect 13287 7295 13313 7321
rect 7575 7239 7601 7265
rect 11327 7239 11353 7265
rect 14631 7239 14657 7265
rect 7967 7183 7993 7209
rect 9815 7127 9841 7153
rect 9871 7155 9897 7181
rect 12895 7127 12921 7153
rect 13063 7127 13089 7153
rect 14743 7127 14769 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8359 6959 8385 6985
rect 11775 6959 11801 6985
rect 8415 6903 8441 6929
rect 10487 6903 10513 6929
rect 10151 6847 10177 6873
rect 11551 6791 11577 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9255 6511 9281 6537
rect 10319 6511 10345 6537
rect 10767 6511 10793 6537
rect 8919 6455 8945 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 12895 2143 12921 2169
rect 13399 2031 13425 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 13063 1807 13089 1833
rect 8807 1751 8833 1777
rect 10375 1751 10401 1777
rect 12615 1751 12641 1777
rect 10879 1639 10905 1665
rect 12279 1639 12305 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 9408 20600 9464 21000
rect 10080 20600 10136 21000
rect 11088 20600 11144 21000
rect 11760 20600 11816 21000
rect 12768 20600 12824 21000
rect 14112 20600 14168 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 9422 19081 9450 20600
rect 9422 19055 9423 19081
rect 9449 19055 9450 19081
rect 9422 19049 9450 19055
rect 9870 19026 9898 19031
rect 9478 19025 9898 19026
rect 9478 18999 9871 19025
rect 9897 18999 9898 19025
rect 9478 18998 9898 18999
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 9478 14042 9506 18998
rect 9870 18993 9898 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10094 18746 10122 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 11774 19138 11802 20600
rect 12782 19306 12810 20600
rect 12782 19273 12810 19278
rect 13398 19306 13426 19311
rect 11774 19105 11802 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 10822 19025 10850 19031
rect 10822 18999 10823 19025
rect 10849 18999 10850 19025
rect 10094 18713 10122 18718
rect 10710 18746 10738 18751
rect 10710 18699 10738 18718
rect 10206 18633 10234 18639
rect 10206 18607 10207 18633
rect 10233 18607 10234 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9814 14209 9842 14215
rect 9814 14183 9815 14209
rect 9841 14183 9842 14209
rect 9478 14041 9674 14042
rect 9478 14015 9479 14041
rect 9505 14015 9674 14041
rect 9478 14014 9674 14015
rect 9478 14009 9506 14014
rect 8974 13985 9002 13991
rect 8974 13959 8975 13985
rect 9001 13959 9002 13985
rect 8862 13930 8890 13935
rect 8582 13929 8890 13930
rect 8582 13903 8863 13929
rect 8889 13903 8890 13929
rect 8582 13902 8890 13903
rect 2086 13818 2114 13823
rect 966 13593 994 13599
rect 966 13567 967 13593
rect 993 13567 994 13593
rect 966 13146 994 13567
rect 966 13113 994 13118
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 966 10738 994 10743
rect 966 10691 994 10710
rect 2086 10290 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8582 13593 8610 13902
rect 8862 13897 8890 13902
rect 8582 13567 8583 13593
rect 8609 13567 8610 13593
rect 8582 13561 8610 13567
rect 2142 13538 2170 13543
rect 2142 13491 2170 13510
rect 6174 13538 6202 13543
rect 6174 13202 6202 13510
rect 8190 13537 8218 13543
rect 8190 13511 8191 13537
rect 8217 13511 8218 13537
rect 7574 13481 7602 13487
rect 7574 13455 7575 13481
rect 7601 13455 7602 13481
rect 7126 13425 7154 13431
rect 7238 13426 7266 13431
rect 7126 13399 7127 13425
rect 7153 13399 7154 13425
rect 7126 13258 7154 13399
rect 7126 13225 7154 13230
rect 7182 13425 7266 13426
rect 7182 13399 7239 13425
rect 7265 13399 7266 13425
rect 7182 13398 7266 13399
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 6062 13146 6090 13151
rect 6062 13089 6090 13118
rect 6062 13063 6063 13089
rect 6089 13063 6090 13089
rect 6062 13057 6090 13063
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6174 12305 6202 13174
rect 7126 13089 7154 13095
rect 7126 13063 7127 13089
rect 7153 13063 7154 13089
rect 7126 12698 7154 13063
rect 7126 12665 7154 12670
rect 6174 12279 6175 12305
rect 6201 12279 6202 12305
rect 6174 12273 6202 12279
rect 7182 12306 7210 13398
rect 7238 13393 7266 13398
rect 7294 13425 7322 13431
rect 7294 13399 7295 13425
rect 7321 13399 7322 13425
rect 7294 12810 7322 13399
rect 7350 13425 7378 13431
rect 7350 13399 7351 13425
rect 7377 13399 7378 13425
rect 7350 12922 7378 13399
rect 7350 12889 7378 12894
rect 7462 13425 7490 13431
rect 7462 13399 7463 13425
rect 7489 13399 7490 13425
rect 7462 12810 7490 13399
rect 7518 13145 7546 13151
rect 7518 13119 7519 13145
rect 7545 13119 7546 13145
rect 7518 12866 7546 13119
rect 7574 13146 7602 13455
rect 7630 13482 7658 13487
rect 7630 13481 7826 13482
rect 7630 13455 7631 13481
rect 7657 13455 7826 13481
rect 7630 13454 7826 13455
rect 7630 13449 7658 13454
rect 7798 13426 7826 13454
rect 7630 13258 7658 13263
rect 7630 13211 7658 13230
rect 7742 13202 7770 13207
rect 7742 13155 7770 13174
rect 7798 13201 7826 13398
rect 7798 13175 7799 13201
rect 7825 13175 7826 13201
rect 7798 13169 7826 13175
rect 7574 13113 7602 13118
rect 8022 13146 8050 13151
rect 8190 13146 8218 13511
rect 8022 13145 8190 13146
rect 8022 13119 8023 13145
rect 8049 13119 8190 13145
rect 8022 13118 8190 13119
rect 8022 13113 8050 13118
rect 8190 13113 8218 13118
rect 8694 13146 8722 13151
rect 7518 12838 7658 12866
rect 7238 12782 7322 12810
rect 7350 12782 7490 12810
rect 7238 12417 7266 12782
rect 7294 12698 7322 12703
rect 7350 12698 7378 12782
rect 7574 12753 7602 12759
rect 7574 12727 7575 12753
rect 7601 12727 7602 12753
rect 7294 12697 7378 12698
rect 7294 12671 7295 12697
rect 7321 12671 7378 12697
rect 7294 12670 7378 12671
rect 7406 12697 7434 12703
rect 7406 12671 7407 12697
rect 7433 12671 7434 12697
rect 7294 12665 7322 12670
rect 7238 12391 7239 12417
rect 7265 12391 7266 12417
rect 7238 12385 7266 12391
rect 7406 12306 7434 12671
rect 7462 12698 7490 12703
rect 7462 12651 7490 12670
rect 7182 12278 7434 12306
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11970 2170 11975
rect 6902 11970 6930 11975
rect 2142 11923 2170 11942
rect 6790 11942 6902 11970
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 6790 11577 6818 11942
rect 6902 11923 6930 11942
rect 6790 11551 6791 11577
rect 6817 11551 6818 11577
rect 5334 11522 5362 11527
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 5334 11018 5362 11494
rect 6398 11521 6426 11527
rect 6398 11495 6399 11521
rect 6425 11495 6426 11521
rect 6398 11130 6426 11495
rect 6398 11097 6426 11102
rect 6622 11186 6650 11191
rect 5334 10985 5362 10990
rect 2142 10794 2170 10799
rect 2142 10747 2170 10766
rect 5222 10794 5250 10799
rect 5222 10737 5250 10766
rect 5222 10711 5223 10737
rect 5249 10711 5250 10737
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 5222 10402 5250 10711
rect 6286 10738 6314 10743
rect 6286 10691 6314 10710
rect 6622 10682 6650 11158
rect 6734 11130 6762 11135
rect 6734 11083 6762 11102
rect 6790 10906 6818 11551
rect 6958 11914 6986 11919
rect 6958 11522 6986 11886
rect 6958 11475 6986 11494
rect 7406 11466 7434 12278
rect 7406 11433 7434 11438
rect 7462 12586 7490 12591
rect 6958 11410 6986 11415
rect 6902 11130 6930 11135
rect 6902 11083 6930 11102
rect 6678 10878 6790 10906
rect 6678 10793 6706 10878
rect 6790 10859 6818 10878
rect 6958 10905 6986 11382
rect 6958 10879 6959 10905
rect 6985 10879 6986 10905
rect 6958 10873 6986 10879
rect 7126 10906 7154 10911
rect 6678 10767 6679 10793
rect 6705 10767 6706 10793
rect 6678 10761 6706 10767
rect 6846 10793 6874 10799
rect 6846 10767 6847 10793
rect 6873 10767 6874 10793
rect 6622 10654 6762 10682
rect 5222 10369 5250 10374
rect 6734 10345 6762 10654
rect 6734 10319 6735 10345
rect 6761 10319 6762 10345
rect 6734 10313 6762 10319
rect 2086 10257 2114 10262
rect 6342 10066 6370 10071
rect 6846 10066 6874 10767
rect 6902 10738 6930 10743
rect 6902 10691 6930 10710
rect 7126 10457 7154 10878
rect 7238 10849 7266 10855
rect 7238 10823 7239 10849
rect 7265 10823 7266 10849
rect 7182 10794 7210 10799
rect 7238 10794 7266 10823
rect 7182 10793 7266 10794
rect 7182 10767 7183 10793
rect 7209 10767 7266 10793
rect 7182 10766 7266 10767
rect 7350 10849 7378 10855
rect 7350 10823 7351 10849
rect 7377 10823 7378 10849
rect 7182 10761 7210 10766
rect 7126 10431 7127 10457
rect 7153 10431 7154 10457
rect 7126 10425 7154 10431
rect 6902 10402 6930 10407
rect 6902 10355 6930 10374
rect 7350 10402 7378 10823
rect 7406 10850 7434 10855
rect 7462 10850 7490 12558
rect 7574 11298 7602 12727
rect 7630 12361 7658 12838
rect 7686 12754 7714 12759
rect 7686 12707 7714 12726
rect 7630 12335 7631 12361
rect 7657 12335 7658 12361
rect 7630 12306 7658 12335
rect 7630 11970 7658 12278
rect 7854 12306 7882 12311
rect 8694 12306 8722 13118
rect 7854 12259 7882 12278
rect 8526 12278 8694 12306
rect 8414 11970 8442 11975
rect 7630 11937 7658 11942
rect 8358 11969 8442 11970
rect 8358 11943 8415 11969
rect 8441 11943 8442 11969
rect 8358 11942 8442 11943
rect 7910 11914 7938 11919
rect 7574 11265 7602 11270
rect 7686 11466 7714 11471
rect 7686 11297 7714 11438
rect 7686 11271 7687 11297
rect 7713 11271 7714 11297
rect 7686 11265 7714 11271
rect 7910 11297 7938 11886
rect 8358 11914 8386 11942
rect 8414 11937 8442 11942
rect 8358 11881 8386 11886
rect 8022 11858 8050 11863
rect 8022 11633 8050 11830
rect 8470 11858 8498 11863
rect 8470 11811 8498 11830
rect 8022 11607 8023 11633
rect 8049 11607 8050 11633
rect 8022 11601 8050 11607
rect 8414 11578 8442 11583
rect 8526 11578 8554 12278
rect 8694 12273 8722 12278
rect 8918 12306 8946 12311
rect 8918 12025 8946 12278
rect 8918 11999 8919 12025
rect 8945 11999 8946 12025
rect 8918 11993 8946 11999
rect 8582 11913 8610 11919
rect 8582 11887 8583 11913
rect 8609 11887 8610 11913
rect 8582 11634 8610 11887
rect 8694 11914 8722 11919
rect 8694 11913 8778 11914
rect 8694 11887 8695 11913
rect 8721 11887 8778 11913
rect 8694 11886 8778 11887
rect 8694 11881 8722 11886
rect 8582 11601 8610 11606
rect 8694 11746 8722 11751
rect 8694 11633 8722 11718
rect 8694 11607 8695 11633
rect 8721 11607 8722 11633
rect 8414 11577 8554 11578
rect 8414 11551 8415 11577
rect 8441 11551 8554 11577
rect 8414 11550 8554 11551
rect 8414 11545 8442 11550
rect 8582 11522 8610 11527
rect 7910 11271 7911 11297
rect 7937 11271 7938 11297
rect 7910 11265 7938 11271
rect 7966 11298 7994 11303
rect 7966 11251 7994 11270
rect 7798 11185 7826 11191
rect 7798 11159 7799 11185
rect 7825 11159 7826 11185
rect 7630 11130 7658 11135
rect 7630 11083 7658 11102
rect 7406 10849 7490 10850
rect 7406 10823 7407 10849
rect 7433 10823 7490 10849
rect 7406 10822 7490 10823
rect 7630 11018 7658 11023
rect 7630 10849 7658 10990
rect 7798 10905 7826 11159
rect 8582 11185 8610 11494
rect 8694 11410 8722 11607
rect 8694 11377 8722 11382
rect 8750 11241 8778 11886
rect 8750 11215 8751 11241
rect 8777 11215 8778 11241
rect 8750 11209 8778 11215
rect 8806 11577 8834 11583
rect 8806 11551 8807 11577
rect 8833 11551 8834 11577
rect 8582 11159 8583 11185
rect 8609 11159 8610 11185
rect 8582 11153 8610 11159
rect 8806 11186 8834 11551
rect 8974 11578 9002 13959
rect 9030 13930 9058 13935
rect 9030 13883 9058 13902
rect 9366 13930 9394 13935
rect 9366 13883 9394 13902
rect 9534 13929 9562 13935
rect 9534 13903 9535 13929
rect 9561 13903 9562 13929
rect 9534 13258 9562 13903
rect 9646 13593 9674 14014
rect 9814 13930 9842 14183
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9870 13930 9898 13935
rect 9814 13902 9870 13930
rect 9870 13883 9898 13902
rect 9870 13650 9898 13655
rect 9646 13567 9647 13593
rect 9673 13567 9674 13593
rect 9646 13561 9674 13567
rect 9702 13649 9898 13650
rect 9702 13623 9871 13649
rect 9897 13623 9898 13649
rect 9702 13622 9898 13623
rect 9702 13454 9730 13622
rect 9870 13617 9898 13622
rect 9870 13538 9898 13543
rect 10206 13538 10234 18607
rect 10262 13873 10290 13879
rect 10262 13847 10263 13873
rect 10289 13847 10290 13873
rect 10262 13650 10290 13847
rect 10822 13874 10850 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 13398 18745 13426 19278
rect 14126 18970 14154 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 14238 18970 14266 18975
rect 14126 18969 14266 18970
rect 14126 18943 14239 18969
rect 14265 18943 14266 18969
rect 14126 18942 14266 18943
rect 14238 18937 14266 18942
rect 13398 18719 13399 18745
rect 13425 18719 13426 18745
rect 13398 18713 13426 18719
rect 12894 18633 12922 18639
rect 12894 18607 12895 18633
rect 12921 18607 12922 18633
rect 12894 15974 12922 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 12110 15946 12306 15974
rect 12670 15946 12922 15974
rect 10318 13650 10346 13655
rect 10262 13649 10346 13650
rect 10262 13623 10319 13649
rect 10345 13623 10346 13649
rect 10262 13622 10346 13623
rect 10318 13617 10346 13622
rect 9534 13225 9562 13230
rect 9646 13426 9730 13454
rect 9814 13481 9842 13487
rect 9814 13455 9815 13481
rect 9841 13455 9842 13481
rect 9814 13426 9842 13455
rect 9870 13481 9898 13510
rect 9870 13455 9871 13481
rect 9897 13455 9898 13481
rect 9870 13449 9898 13455
rect 10150 13510 10206 13538
rect 9086 13090 9114 13095
rect 9086 13089 9394 13090
rect 9086 13063 9087 13089
rect 9113 13063 9394 13089
rect 9086 13062 9394 13063
rect 9086 13057 9114 13062
rect 9366 12809 9394 13062
rect 9366 12783 9367 12809
rect 9393 12783 9394 12809
rect 9366 12777 9394 12783
rect 9086 12754 9114 12759
rect 8862 11466 8890 11471
rect 8862 11419 8890 11438
rect 8974 11242 9002 11550
rect 8806 11153 8834 11158
rect 8918 11214 9002 11242
rect 9030 11634 9058 11639
rect 8694 11074 8722 11079
rect 8806 11074 8834 11079
rect 8694 11073 8806 11074
rect 8694 11047 8695 11073
rect 8721 11047 8806 11073
rect 8694 11046 8806 11047
rect 8694 11041 8722 11046
rect 8806 11041 8834 11046
rect 8862 11073 8890 11079
rect 8862 11047 8863 11073
rect 8889 11047 8890 11073
rect 8862 10962 8890 11047
rect 7798 10879 7799 10905
rect 7825 10879 7826 10905
rect 7798 10873 7826 10879
rect 8694 10934 8890 10962
rect 7630 10823 7631 10849
rect 7657 10823 7658 10849
rect 7406 10817 7434 10822
rect 7630 10817 7658 10823
rect 7350 10369 7378 10374
rect 7742 10793 7770 10799
rect 7742 10767 7743 10793
rect 7769 10767 7770 10793
rect 6342 10019 6370 10038
rect 6734 10038 6846 10066
rect 6006 10009 6034 10015
rect 6006 9983 6007 10009
rect 6033 9983 6034 10009
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 6006 9226 6034 9983
rect 6734 9561 6762 10038
rect 6846 10033 6874 10038
rect 7406 10010 7434 10015
rect 7406 9953 7434 9982
rect 7406 9927 7407 9953
rect 7433 9927 7434 9953
rect 7406 9921 7434 9927
rect 7686 9953 7714 9959
rect 7686 9927 7687 9953
rect 7713 9927 7714 9953
rect 6902 9898 6930 9903
rect 6902 9617 6930 9870
rect 6902 9591 6903 9617
rect 6929 9591 6930 9617
rect 6902 9585 6930 9591
rect 6734 9535 6735 9561
rect 6761 9535 6762 9561
rect 6734 9529 6762 9535
rect 7294 9506 7322 9511
rect 6006 9193 6034 9198
rect 7014 9225 7042 9231
rect 7014 9199 7015 9225
rect 7041 9199 7042 9225
rect 6398 9170 6426 9175
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5614 8834 5642 8839
rect 2142 8441 2170 8447
rect 2142 8415 2143 8441
rect 2169 8415 2170 8441
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 966 8073 994 8078
rect 2142 7602 2170 8415
rect 5614 8385 5642 8806
rect 5614 8359 5615 8385
rect 5641 8359 5642 8385
rect 5614 8353 5642 8359
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6398 8105 6426 9142
rect 7014 8554 7042 9199
rect 7182 9225 7210 9231
rect 7182 9199 7183 9225
rect 7209 9199 7210 9225
rect 7126 9170 7154 9175
rect 7126 9123 7154 9142
rect 7182 8834 7210 9199
rect 7182 8801 7210 8806
rect 6902 8526 7042 8554
rect 7294 8553 7322 9478
rect 7350 9225 7378 9231
rect 7350 9199 7351 9225
rect 7377 9199 7378 9225
rect 7350 9058 7378 9199
rect 7518 9226 7546 9231
rect 7686 9226 7714 9927
rect 7742 9506 7770 10767
rect 7854 10793 7882 10799
rect 7854 10767 7855 10793
rect 7881 10767 7882 10793
rect 7854 10122 7882 10767
rect 7966 10794 7994 10799
rect 7966 10747 7994 10766
rect 7854 10089 7882 10094
rect 8022 10458 8050 10463
rect 8022 10065 8050 10430
rect 8638 10458 8666 10463
rect 8638 10411 8666 10430
rect 8526 10122 8554 10127
rect 8694 10122 8722 10934
rect 8918 10905 8946 11214
rect 9030 11186 9058 11606
rect 8918 10879 8919 10905
rect 8945 10879 8946 10905
rect 8918 10873 8946 10879
rect 8974 11130 9002 11135
rect 8806 10850 8834 10855
rect 8806 10849 8890 10850
rect 8806 10823 8807 10849
rect 8833 10823 8890 10849
rect 8806 10822 8890 10823
rect 8806 10817 8834 10822
rect 8750 10794 8778 10799
rect 8750 10747 8778 10766
rect 8806 10402 8834 10407
rect 8862 10402 8890 10822
rect 8806 10401 8890 10402
rect 8806 10375 8807 10401
rect 8833 10375 8890 10401
rect 8806 10374 8890 10375
rect 8694 10094 8778 10122
rect 8022 10039 8023 10065
rect 8049 10039 8050 10065
rect 8022 10033 8050 10039
rect 8358 10065 8386 10071
rect 8358 10039 8359 10065
rect 8385 10039 8386 10065
rect 8246 10009 8274 10015
rect 8246 9983 8247 10009
rect 8273 9983 8274 10009
rect 7966 9898 7994 9903
rect 7966 9851 7994 9870
rect 8134 9898 8162 9903
rect 8134 9851 8162 9870
rect 7742 9473 7770 9478
rect 8246 9506 8274 9983
rect 8358 9898 8386 10039
rect 8470 10066 8498 10071
rect 8414 10009 8442 10015
rect 8414 9983 8415 10009
rect 8441 9983 8442 10009
rect 8414 9954 8442 9983
rect 8414 9921 8442 9926
rect 8358 9730 8386 9870
rect 8414 9730 8442 9735
rect 8358 9729 8442 9730
rect 8358 9703 8415 9729
rect 8441 9703 8442 9729
rect 8358 9702 8442 9703
rect 8414 9697 8442 9702
rect 8470 9561 8498 10038
rect 8470 9535 8471 9561
rect 8497 9535 8498 9561
rect 8470 9529 8498 9535
rect 8246 9473 8274 9478
rect 8526 9450 8554 10094
rect 8694 10010 8722 10015
rect 8694 9963 8722 9982
rect 8750 9842 8778 10094
rect 8750 9809 8778 9814
rect 8750 9730 8778 9735
rect 8806 9730 8834 10374
rect 8862 10066 8890 10071
rect 8862 10065 8946 10066
rect 8862 10039 8863 10065
rect 8889 10039 8946 10065
rect 8862 10038 8946 10039
rect 8862 10033 8890 10038
rect 8750 9729 8834 9730
rect 8750 9703 8751 9729
rect 8777 9703 8834 9729
rect 8750 9702 8834 9703
rect 8862 9842 8890 9847
rect 8750 9697 8778 9702
rect 7546 9198 7714 9226
rect 8470 9422 8554 9450
rect 8582 9561 8610 9567
rect 8582 9535 8583 9561
rect 8609 9535 8610 9561
rect 7518 9193 7546 9198
rect 7350 9025 7378 9030
rect 7294 8527 7295 8553
rect 7321 8527 7322 8553
rect 6678 8386 6706 8391
rect 6454 8385 6706 8386
rect 6454 8359 6679 8385
rect 6705 8359 6706 8385
rect 6454 8358 6706 8359
rect 6454 8161 6482 8358
rect 6678 8353 6706 8358
rect 6454 8135 6455 8161
rect 6481 8135 6482 8161
rect 6454 8129 6482 8135
rect 6398 8079 6399 8105
rect 6425 8079 6426 8105
rect 6398 8073 6426 8079
rect 6902 8050 6930 8526
rect 7294 8521 7322 8527
rect 7574 8553 7602 9198
rect 7574 8527 7575 8553
rect 7601 8527 7602 8553
rect 7014 8441 7042 8447
rect 7238 8442 7266 8447
rect 7014 8415 7015 8441
rect 7041 8415 7042 8441
rect 7014 8386 7042 8415
rect 7014 8353 7042 8358
rect 7070 8441 7266 8442
rect 7070 8415 7239 8441
rect 7265 8415 7266 8441
rect 7070 8414 7266 8415
rect 7070 8218 7098 8414
rect 7238 8409 7266 8414
rect 7574 8386 7602 8527
rect 7294 8330 7322 8335
rect 6958 8190 7098 8218
rect 7126 8329 7322 8330
rect 7126 8303 7295 8329
rect 7321 8303 7322 8329
rect 7126 8302 7322 8303
rect 6958 8161 6986 8190
rect 6958 8135 6959 8161
rect 6985 8135 6986 8161
rect 6958 8129 6986 8135
rect 6902 8022 7042 8050
rect 7014 7993 7042 8022
rect 7014 7967 7015 7993
rect 7041 7967 7042 7993
rect 6958 7938 6986 7943
rect 6902 7937 6986 7938
rect 6902 7911 6959 7937
rect 6985 7911 6986 7937
rect 6902 7910 6986 7911
rect 2142 7569 2170 7574
rect 5894 7602 5922 7607
rect 5894 7555 5922 7574
rect 6846 7602 6874 7607
rect 6902 7602 6930 7910
rect 6958 7905 6986 7910
rect 7014 7938 7042 7967
rect 7014 7905 7042 7910
rect 7126 7826 7154 8302
rect 7294 8297 7322 8302
rect 6958 7798 7154 7826
rect 7574 8049 7602 8358
rect 7910 8722 7938 8727
rect 7910 8105 7938 8694
rect 8358 8722 8386 8727
rect 8470 8722 8498 9422
rect 8582 9338 8610 9535
rect 8582 9305 8610 9310
rect 8526 8834 8554 8839
rect 8806 8834 8834 8839
rect 8526 8833 8834 8834
rect 8526 8807 8527 8833
rect 8553 8807 8807 8833
rect 8833 8807 8834 8833
rect 8526 8806 8834 8807
rect 8526 8801 8554 8806
rect 8750 8722 8778 8727
rect 8470 8721 8778 8722
rect 8470 8695 8751 8721
rect 8777 8695 8778 8721
rect 8470 8694 8778 8695
rect 8358 8675 8386 8694
rect 8750 8330 8778 8694
rect 8806 8553 8834 8806
rect 8862 8666 8890 9814
rect 8918 9617 8946 10038
rect 8918 9591 8919 9617
rect 8945 9591 8946 9617
rect 8918 9506 8946 9591
rect 8974 9506 9002 11102
rect 9030 10906 9058 11158
rect 9086 11074 9114 12726
rect 9254 12754 9282 12759
rect 9254 12473 9282 12726
rect 9646 12753 9674 13426
rect 9646 12727 9647 12753
rect 9673 12727 9674 12753
rect 9646 12721 9674 12727
rect 9814 12754 9842 13398
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9814 12707 9842 12726
rect 9926 13258 9954 13263
rect 9926 12697 9954 13230
rect 10150 13089 10178 13510
rect 10206 13505 10234 13510
rect 10374 13482 10402 13487
rect 10710 13482 10738 13487
rect 10374 13481 10738 13482
rect 10374 13455 10375 13481
rect 10401 13455 10711 13481
rect 10737 13455 10738 13481
rect 10374 13454 10738 13455
rect 10374 13449 10402 13454
rect 10710 13449 10738 13454
rect 10822 13481 10850 13846
rect 11326 13874 11354 13879
rect 11326 13827 11354 13846
rect 11550 13873 11578 13879
rect 11550 13847 11551 13873
rect 11577 13847 11578 13873
rect 10822 13455 10823 13481
rect 10849 13455 10850 13481
rect 10822 13449 10850 13455
rect 10878 13482 10906 13487
rect 11550 13454 11578 13847
rect 12110 13454 12138 15946
rect 10878 13435 10906 13454
rect 10150 13063 10151 13089
rect 10177 13063 10178 13089
rect 10150 13057 10178 13063
rect 10318 13425 10346 13431
rect 10318 13399 10319 13425
rect 10345 13399 10346 13425
rect 9926 12671 9927 12697
rect 9953 12671 9954 12697
rect 9926 12665 9954 12671
rect 9310 12642 9338 12647
rect 9422 12642 9450 12647
rect 9310 12641 9394 12642
rect 9310 12615 9311 12641
rect 9337 12615 9394 12641
rect 9310 12614 9394 12615
rect 9310 12609 9338 12614
rect 9254 12447 9255 12473
rect 9281 12447 9282 12473
rect 9254 12441 9282 12447
rect 9310 11578 9338 11583
rect 9310 11531 9338 11550
rect 9198 11354 9226 11359
rect 9198 11185 9226 11326
rect 9198 11159 9199 11185
rect 9225 11159 9226 11185
rect 9198 11153 9226 11159
rect 9086 11027 9114 11046
rect 9086 10906 9114 10911
rect 9030 10905 9114 10906
rect 9030 10879 9087 10905
rect 9113 10879 9114 10905
rect 9030 10878 9114 10879
rect 9086 10873 9114 10878
rect 9198 10850 9226 10855
rect 9142 10794 9170 10799
rect 9086 10402 9114 10407
rect 9086 10355 9114 10374
rect 9030 10345 9058 10351
rect 9030 10319 9031 10345
rect 9057 10319 9058 10345
rect 9030 10010 9058 10319
rect 9030 9977 9058 9982
rect 9142 10010 9170 10766
rect 9198 10793 9226 10822
rect 9198 10767 9199 10793
rect 9225 10767 9226 10793
rect 9198 10066 9226 10767
rect 9198 10019 9226 10038
rect 9142 9977 9170 9982
rect 9310 9897 9338 9903
rect 9310 9871 9311 9897
rect 9337 9871 9338 9897
rect 9030 9618 9058 9623
rect 9254 9618 9282 9623
rect 9030 9617 9282 9618
rect 9030 9591 9031 9617
rect 9057 9591 9255 9617
rect 9281 9591 9282 9617
rect 9030 9590 9282 9591
rect 9030 9585 9058 9590
rect 8974 9478 9058 9506
rect 8918 9473 8946 9478
rect 8974 9338 9002 9343
rect 8918 9226 8946 9231
rect 8974 9226 9002 9310
rect 8918 9225 9002 9226
rect 8918 9199 8919 9225
rect 8945 9199 9002 9225
rect 8918 9198 9002 9199
rect 8918 9193 8946 9198
rect 8974 8889 9002 9198
rect 9030 9337 9058 9478
rect 9030 9311 9031 9337
rect 9057 9311 9058 9337
rect 9030 9226 9058 9311
rect 9030 9193 9058 9198
rect 8974 8863 8975 8889
rect 9001 8863 9002 8889
rect 8974 8857 9002 8863
rect 8862 8633 8890 8638
rect 9086 8554 9114 9590
rect 9254 9562 9282 9590
rect 9254 9529 9282 9534
rect 9310 9506 9338 9871
rect 9310 9473 9338 9478
rect 9310 9338 9338 9343
rect 9366 9338 9394 12614
rect 9422 12641 9674 12642
rect 9422 12615 9423 12641
rect 9449 12615 9674 12641
rect 9422 12614 9674 12615
rect 9422 12609 9450 12614
rect 9422 12362 9450 12367
rect 9422 12361 9506 12362
rect 9422 12335 9423 12361
rect 9449 12335 9506 12361
rect 9422 12334 9506 12335
rect 9422 12329 9450 12334
rect 9478 10402 9506 12334
rect 9590 11690 9618 11695
rect 9534 11578 9562 11583
rect 9590 11578 9618 11662
rect 9646 11634 9674 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9646 11601 9674 11606
rect 9814 12361 9842 12367
rect 9814 12335 9815 12361
rect 9841 12335 9842 12361
rect 9534 11577 9618 11578
rect 9534 11551 9535 11577
rect 9561 11551 9618 11577
rect 9534 11550 9618 11551
rect 9534 11545 9562 11550
rect 9590 10849 9618 11550
rect 9758 11465 9786 11471
rect 9758 11439 9759 11465
rect 9785 11439 9786 11465
rect 9758 11298 9786 11439
rect 9758 11265 9786 11270
rect 9590 10823 9591 10849
rect 9617 10823 9618 10849
rect 9590 10817 9618 10823
rect 9702 10794 9730 10813
rect 9702 10761 9730 10766
rect 9646 10458 9674 10463
rect 9590 10430 9646 10458
rect 9478 10374 9562 10402
rect 9478 10290 9506 10295
rect 9478 10243 9506 10262
rect 9422 10066 9450 10071
rect 9422 9673 9450 10038
rect 9478 9898 9506 9903
rect 9478 9851 9506 9870
rect 9422 9647 9423 9673
rect 9449 9647 9450 9673
rect 9422 9641 9450 9647
rect 9310 9337 9394 9338
rect 9310 9311 9311 9337
rect 9337 9311 9394 9337
rect 9310 9310 9394 9311
rect 9310 9305 9338 9310
rect 9142 9226 9170 9231
rect 9142 9179 9170 9198
rect 9310 9225 9338 9231
rect 9310 9199 9311 9225
rect 9337 9199 9338 9225
rect 9310 8722 9338 9199
rect 9366 9226 9394 9231
rect 9366 8833 9394 9198
rect 9478 9225 9506 9231
rect 9478 9199 9479 9225
rect 9505 9199 9506 9225
rect 9478 8889 9506 9199
rect 9534 9226 9562 10374
rect 9534 9193 9562 9198
rect 9478 8863 9479 8889
rect 9505 8863 9506 8889
rect 9478 8857 9506 8863
rect 9366 8807 9367 8833
rect 9393 8807 9394 8833
rect 9366 8801 9394 8807
rect 9590 8834 9618 10430
rect 9646 10425 9674 10430
rect 9646 10290 9674 10295
rect 9646 10009 9674 10262
rect 9814 10066 9842 12335
rect 10038 11969 10066 11975
rect 10038 11943 10039 11969
rect 10065 11943 10066 11969
rect 9870 11913 9898 11919
rect 9870 11887 9871 11913
rect 9897 11887 9898 11913
rect 9870 11858 9898 11887
rect 9926 11914 9954 11919
rect 9926 11867 9954 11886
rect 10038 11858 10066 11943
rect 10038 11830 10122 11858
rect 9870 11825 9898 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11578 10122 11830
rect 10318 11690 10346 13399
rect 11494 13426 11578 13454
rect 11998 13426 12026 13431
rect 10374 13314 10402 13319
rect 10374 13089 10402 13286
rect 10374 13063 10375 13089
rect 10401 13063 10402 13089
rect 10374 12306 10402 13063
rect 11494 12753 11522 13426
rect 11494 12727 11495 12753
rect 11521 12727 11522 12753
rect 11270 12642 11298 12647
rect 11494 12642 11522 12727
rect 11270 12641 11522 12642
rect 11270 12615 11271 12641
rect 11297 12615 11522 12641
rect 11270 12614 11522 12615
rect 11270 12609 11298 12614
rect 10374 12273 10402 12278
rect 10710 12306 10738 12311
rect 10710 11969 10738 12278
rect 11494 12306 11522 12614
rect 11494 12273 11522 12278
rect 11550 13146 11578 13151
rect 11550 12642 11578 13118
rect 11550 12194 11578 12614
rect 10710 11943 10711 11969
rect 10737 11943 10738 11969
rect 10710 11937 10738 11943
rect 11438 12166 11578 12194
rect 11662 13145 11690 13151
rect 11662 13119 11663 13145
rect 11689 13119 11690 13145
rect 10318 11657 10346 11662
rect 10990 11914 11018 11919
rect 10206 11578 10234 11583
rect 10094 11550 10206 11578
rect 10038 11522 10066 11527
rect 10038 11475 10066 11494
rect 9926 11466 9954 11471
rect 9926 11465 10010 11466
rect 9926 11439 9927 11465
rect 9953 11439 10010 11465
rect 9926 11438 10010 11439
rect 9926 11433 9954 11438
rect 9982 11242 10010 11438
rect 10150 11242 10178 11247
rect 9982 11214 10150 11242
rect 10150 11195 10178 11214
rect 10094 11130 10122 11135
rect 10206 11130 10234 11550
rect 10318 11577 10346 11583
rect 10318 11551 10319 11577
rect 10345 11551 10346 11577
rect 10262 11522 10290 11527
rect 10262 11475 10290 11494
rect 10318 11410 10346 11551
rect 10262 11186 10290 11191
rect 10318 11186 10346 11382
rect 10290 11158 10346 11186
rect 10542 11577 10570 11583
rect 10542 11551 10543 11577
rect 10569 11551 10570 11577
rect 10262 11139 10290 11158
rect 10094 11129 10234 11130
rect 10094 11103 10095 11129
rect 10121 11103 10234 11129
rect 10094 11102 10234 11103
rect 10374 11130 10402 11135
rect 10374 11129 10514 11130
rect 10374 11103 10375 11129
rect 10401 11103 10514 11129
rect 10374 11102 10514 11103
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10094 10906 10122 11102
rect 10374 11097 10402 11102
rect 10038 10878 10122 10906
rect 9870 10794 9898 10799
rect 9870 10402 9898 10766
rect 9870 10355 9898 10374
rect 10038 10345 10066 10878
rect 10374 10850 10402 10855
rect 10374 10803 10402 10822
rect 10038 10319 10039 10345
rect 10065 10319 10066 10345
rect 10038 10313 10066 10319
rect 10318 10402 10346 10407
rect 10486 10402 10514 11102
rect 10542 10906 10570 11551
rect 10598 11578 10626 11583
rect 10598 11531 10626 11550
rect 10766 11577 10794 11583
rect 10766 11551 10767 11577
rect 10793 11551 10794 11577
rect 10710 11354 10738 11359
rect 10654 11242 10682 11247
rect 10654 11185 10682 11214
rect 10654 11159 10655 11185
rect 10681 11159 10682 11185
rect 10654 11153 10682 11159
rect 10542 10873 10570 10878
rect 10598 10402 10626 10407
rect 10486 10401 10626 10402
rect 10486 10375 10599 10401
rect 10625 10375 10626 10401
rect 10486 10374 10626 10375
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9646 9983 9647 10009
rect 9673 9983 9674 10009
rect 9646 9977 9674 9983
rect 9702 10038 9814 10066
rect 9646 9506 9674 9511
rect 9646 9282 9674 9478
rect 9646 9249 9674 9254
rect 9590 8801 9618 8806
rect 9310 8689 9338 8694
rect 9534 8777 9562 8783
rect 9534 8751 9535 8777
rect 9561 8751 9562 8777
rect 9534 8722 9562 8751
rect 9534 8689 9562 8694
rect 8806 8527 8807 8553
rect 8833 8527 8834 8553
rect 8806 8521 8834 8527
rect 8862 8526 9114 8554
rect 8862 8497 8890 8526
rect 8862 8471 8863 8497
rect 8889 8471 8890 8497
rect 8862 8465 8890 8471
rect 8750 8297 8778 8302
rect 8918 8442 8946 8447
rect 7910 8079 7911 8105
rect 7937 8079 7938 8105
rect 7910 8073 7938 8079
rect 7574 8023 7575 8049
rect 7601 8023 7602 8049
rect 6958 7713 6986 7798
rect 7574 7770 7602 8023
rect 6958 7687 6959 7713
rect 6985 7687 6986 7713
rect 6958 7681 6986 7687
rect 7350 7769 7602 7770
rect 7350 7743 7575 7769
rect 7601 7743 7602 7769
rect 7350 7742 7602 7743
rect 7350 7657 7378 7742
rect 7350 7631 7351 7657
rect 7377 7631 7378 7657
rect 7350 7625 7378 7631
rect 6874 7574 6930 7602
rect 7574 7602 7602 7742
rect 6846 7569 6874 7574
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7574 7265 7602 7574
rect 7574 7239 7575 7265
rect 7601 7239 7602 7265
rect 7574 7233 7602 7239
rect 8414 7742 8890 7770
rect 7966 7210 7994 7215
rect 7966 7209 8386 7210
rect 7966 7183 7967 7209
rect 7993 7183 8386 7209
rect 7966 7182 8386 7183
rect 7966 7177 7994 7182
rect 8358 6985 8386 7182
rect 8358 6959 8359 6985
rect 8385 6959 8386 6985
rect 8358 6953 8386 6959
rect 8414 6929 8442 7742
rect 8862 7713 8890 7742
rect 8918 7769 8946 8414
rect 8974 8105 9002 8526
rect 9702 8441 9730 10038
rect 9814 10033 9842 10038
rect 10262 9842 10290 9847
rect 10206 9730 10234 9735
rect 10206 9683 10234 9702
rect 10262 9673 10290 9814
rect 10262 9647 10263 9673
rect 10289 9647 10290 9673
rect 10262 9641 10290 9647
rect 10150 9562 10178 9567
rect 9814 9505 9842 9511
rect 9814 9479 9815 9505
rect 9841 9479 9842 9505
rect 9814 9338 9842 9479
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9814 9305 9842 9310
rect 10150 9337 10178 9534
rect 10318 9561 10346 10374
rect 10598 9786 10626 10374
rect 10598 9753 10626 9758
rect 10710 9673 10738 11326
rect 10710 9647 10711 9673
rect 10737 9647 10738 9673
rect 10710 9641 10738 9647
rect 10598 9618 10626 9623
rect 10318 9535 10319 9561
rect 10345 9535 10346 9561
rect 10318 9529 10346 9535
rect 10374 9617 10626 9618
rect 10374 9591 10599 9617
rect 10625 9591 10626 9617
rect 10374 9590 10626 9591
rect 10262 9338 10290 9343
rect 10374 9338 10402 9590
rect 10598 9585 10626 9590
rect 10766 9394 10794 11551
rect 10990 11577 11018 11886
rect 11046 11913 11074 11919
rect 11046 11887 11047 11913
rect 11073 11887 11074 11913
rect 11046 11689 11074 11887
rect 11046 11663 11047 11689
rect 11073 11663 11074 11689
rect 11046 11657 11074 11663
rect 10990 11551 10991 11577
rect 11017 11551 11018 11577
rect 10990 11545 11018 11551
rect 11046 11578 11074 11583
rect 10878 11466 10906 11471
rect 10878 11419 10906 11438
rect 10934 10849 10962 10855
rect 10934 10823 10935 10849
rect 10961 10823 10962 10849
rect 10934 10570 10962 10823
rect 10878 10542 10934 10570
rect 10878 9730 10906 10542
rect 10934 10537 10962 10542
rect 10990 10402 11018 10407
rect 10990 10355 11018 10374
rect 10934 10066 10962 10071
rect 10934 10019 10962 10038
rect 10878 9617 10906 9702
rect 10878 9591 10879 9617
rect 10905 9591 10906 9617
rect 10150 9311 10151 9337
rect 10177 9311 10178 9337
rect 10150 9305 10178 9311
rect 10206 9337 10402 9338
rect 10206 9311 10263 9337
rect 10289 9311 10402 9337
rect 10206 9310 10402 9311
rect 10430 9366 10794 9394
rect 10822 9561 10850 9567
rect 10822 9535 10823 9561
rect 10849 9535 10850 9561
rect 9702 8415 9703 8441
rect 9729 8415 9730 8441
rect 9702 8409 9730 8415
rect 9758 9281 9786 9287
rect 9758 9255 9759 9281
rect 9785 9255 9786 9281
rect 8974 8079 8975 8105
rect 9001 8079 9002 8105
rect 8974 8073 9002 8079
rect 9030 8330 9058 8335
rect 8918 7743 8919 7769
rect 8945 7743 8946 7769
rect 8918 7737 8946 7743
rect 8862 7687 8863 7713
rect 8889 7687 8890 7713
rect 8862 7681 8890 7687
rect 9030 7713 9058 8302
rect 9030 7687 9031 7713
rect 9057 7687 9058 7713
rect 9030 7681 9058 7687
rect 9198 7937 9226 7943
rect 9198 7911 9199 7937
rect 9225 7911 9226 7937
rect 8750 7658 8778 7663
rect 8750 7611 8778 7630
rect 8806 7657 8834 7663
rect 8806 7631 8807 7657
rect 8833 7631 8834 7657
rect 8806 7490 8834 7631
rect 9198 7602 9226 7911
rect 9758 7658 9786 9255
rect 10094 9282 10122 9287
rect 10094 9235 10122 9254
rect 9870 9226 9898 9231
rect 9870 9179 9898 9198
rect 9814 8834 9842 8839
rect 9814 8787 9842 8806
rect 9870 8722 9898 8741
rect 9870 8689 9898 8694
rect 9982 8722 10010 8727
rect 10150 8722 10178 8727
rect 9982 8721 10122 8722
rect 9982 8695 9983 8721
rect 10009 8695 10122 8721
rect 9982 8694 10122 8695
rect 9982 8689 10010 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10094 8050 10122 8694
rect 10150 8675 10178 8694
rect 10206 8050 10234 9310
rect 10262 9305 10290 9310
rect 10430 9282 10458 9366
rect 10822 9338 10850 9535
rect 10822 9305 10850 9310
rect 10318 9254 10458 9282
rect 10654 9282 10682 9287
rect 10318 8889 10346 9254
rect 10318 8863 10319 8889
rect 10345 8863 10346 8889
rect 10318 8857 10346 8863
rect 10654 8833 10682 9254
rect 10878 9169 10906 9591
rect 11046 9562 11074 11550
rect 11102 11577 11130 11583
rect 11102 11551 11103 11577
rect 11129 11551 11130 11577
rect 11102 11410 11130 11551
rect 11102 11377 11130 11382
rect 11158 11522 11186 11527
rect 11158 11185 11186 11494
rect 11438 11465 11466 12166
rect 11606 11746 11634 11751
rect 11606 11577 11634 11718
rect 11606 11551 11607 11577
rect 11633 11551 11634 11577
rect 11606 11545 11634 11551
rect 11438 11439 11439 11465
rect 11465 11439 11466 11465
rect 11438 11410 11466 11439
rect 11494 11521 11522 11527
rect 11494 11495 11495 11521
rect 11521 11495 11522 11521
rect 11494 11466 11522 11495
rect 11494 11433 11522 11438
rect 11158 11159 11159 11185
rect 11185 11159 11186 11185
rect 11158 11153 11186 11159
rect 11270 11382 11466 11410
rect 11270 11074 11298 11382
rect 11662 11241 11690 13119
rect 11774 13146 11802 13151
rect 11774 13099 11802 13118
rect 11886 13146 11914 13151
rect 11886 13099 11914 13118
rect 11998 13145 12026 13398
rect 11998 13119 11999 13145
rect 12025 13119 12026 13145
rect 11830 13089 11858 13095
rect 11830 13063 11831 13089
rect 11857 13063 11858 13089
rect 11830 12809 11858 13063
rect 11830 12783 11831 12809
rect 11857 12783 11858 12809
rect 11830 12777 11858 12783
rect 11998 11858 12026 13119
rect 11998 11825 12026 11830
rect 12054 13426 12138 13454
rect 12054 12026 12082 13426
rect 12670 13202 12698 15946
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12670 13201 12922 13202
rect 12670 13175 12671 13201
rect 12697 13175 12922 13201
rect 12670 13174 12922 13175
rect 12670 13169 12698 13174
rect 12614 13146 12642 13151
rect 12614 13099 12642 13118
rect 12894 12809 12922 13174
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 12894 12783 12895 12809
rect 12921 12783 12922 12809
rect 12894 12777 12922 12783
rect 13286 12753 13314 12759
rect 13286 12727 13287 12753
rect 13313 12727 13314 12753
rect 13118 12641 13146 12647
rect 13118 12615 13119 12641
rect 13145 12615 13146 12641
rect 13006 12362 13034 12367
rect 13118 12362 13146 12615
rect 13286 12642 13314 12727
rect 13454 12698 13482 12703
rect 13454 12697 13986 12698
rect 13454 12671 13455 12697
rect 13481 12671 13986 12697
rect 13454 12670 13986 12671
rect 13454 12665 13482 12670
rect 13286 12609 13314 12614
rect 13398 12641 13426 12647
rect 13398 12615 13399 12641
rect 13425 12615 13426 12641
rect 13398 12417 13426 12615
rect 13398 12391 13399 12417
rect 13425 12391 13426 12417
rect 13398 12385 13426 12391
rect 13006 12361 13146 12362
rect 13006 12335 13007 12361
rect 13033 12335 13146 12361
rect 13006 12334 13146 12335
rect 12110 12306 12138 12311
rect 12166 12306 12194 12311
rect 12110 12305 12166 12306
rect 12110 12279 12111 12305
rect 12137 12279 12166 12305
rect 12110 12278 12166 12279
rect 12110 12273 12138 12278
rect 12110 12026 12138 12031
rect 12054 12025 12138 12026
rect 12054 11999 12111 12025
rect 12137 11999 12138 12025
rect 12054 11998 12138 11999
rect 12054 11746 12082 11998
rect 12110 11993 12138 11998
rect 12166 11970 12194 12278
rect 12670 12306 12698 12311
rect 12670 12259 12698 12278
rect 13006 12306 13034 12334
rect 13006 12273 13034 12278
rect 13734 12026 13762 12031
rect 12278 11970 12306 11975
rect 12166 11969 12306 11970
rect 12166 11943 12279 11969
rect 12305 11943 12306 11969
rect 12166 11942 12306 11943
rect 12054 11713 12082 11718
rect 11830 11634 11858 11639
rect 11830 11577 11858 11606
rect 12054 11634 12082 11639
rect 12054 11587 12082 11606
rect 11830 11551 11831 11577
rect 11857 11551 11858 11577
rect 11830 11545 11858 11551
rect 12166 11577 12194 11583
rect 12166 11551 12167 11577
rect 12193 11551 12194 11577
rect 11886 11466 11914 11471
rect 11886 11465 11970 11466
rect 11886 11439 11887 11465
rect 11913 11439 11970 11465
rect 11886 11438 11970 11439
rect 11886 11433 11914 11438
rect 11662 11215 11663 11241
rect 11689 11215 11690 11241
rect 11662 11209 11690 11215
rect 11606 11185 11634 11191
rect 11606 11159 11607 11185
rect 11633 11159 11634 11185
rect 11326 11130 11354 11135
rect 11326 11129 11466 11130
rect 11326 11103 11327 11129
rect 11353 11103 11466 11129
rect 11326 11102 11466 11103
rect 11326 11097 11354 11102
rect 11158 11046 11298 11074
rect 11158 10513 11186 11046
rect 11270 10793 11298 10799
rect 11270 10767 11271 10793
rect 11297 10767 11298 10793
rect 11158 10487 11159 10513
rect 11185 10487 11186 10513
rect 11158 10481 11186 10487
rect 11214 10738 11242 10743
rect 11214 10458 11242 10710
rect 11214 10411 11242 10430
rect 11102 9786 11130 9791
rect 11130 9758 11186 9786
rect 11102 9753 11130 9758
rect 10878 9143 10879 9169
rect 10905 9143 10906 9169
rect 10878 9137 10906 9143
rect 10934 9534 11074 9562
rect 10654 8807 10655 8833
rect 10681 8807 10682 8833
rect 10654 8801 10682 8807
rect 10262 8778 10290 8783
rect 10262 8731 10290 8750
rect 10710 8778 10738 8783
rect 10710 8731 10738 8750
rect 10374 8721 10402 8727
rect 10374 8695 10375 8721
rect 10401 8695 10402 8721
rect 10262 8050 10290 8055
rect 10206 8049 10290 8050
rect 10206 8023 10263 8049
rect 10289 8023 10290 8049
rect 10206 8022 10290 8023
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9926 7770 9954 7775
rect 9926 7723 9954 7742
rect 10038 7770 10066 7775
rect 10094 7770 10122 8022
rect 10262 8017 10290 8022
rect 10318 7994 10346 7999
rect 10374 7994 10402 8695
rect 10934 8386 10962 9534
rect 11158 9282 11186 9758
rect 11270 9618 11298 10767
rect 11438 10289 11466 11102
rect 11550 11129 11578 11135
rect 11550 11103 11551 11129
rect 11577 11103 11578 11129
rect 11494 10738 11522 10743
rect 11494 10691 11522 10710
rect 11550 10458 11578 11103
rect 11606 10682 11634 11159
rect 11942 10850 11970 11438
rect 12166 11186 12194 11551
rect 11942 10803 11970 10822
rect 12054 11158 12194 11186
rect 11718 10793 11746 10799
rect 11718 10767 11719 10793
rect 11745 10767 11746 10793
rect 11606 10654 11690 10682
rect 11438 10263 11439 10289
rect 11465 10263 11466 10289
rect 11326 9618 11354 9623
rect 11270 9590 11326 9618
rect 11326 9571 11354 9590
rect 11438 9394 11466 10263
rect 11494 10430 11578 10458
rect 11606 10570 11634 10575
rect 11494 10010 11522 10430
rect 11606 10401 11634 10542
rect 11606 10375 11607 10401
rect 11633 10375 11634 10401
rect 11606 10369 11634 10375
rect 11662 10122 11690 10654
rect 11718 10402 11746 10767
rect 11886 10458 11914 10463
rect 12054 10458 12082 11158
rect 12110 11074 12138 11079
rect 12110 11073 12194 11074
rect 12110 11047 12111 11073
rect 12137 11047 12194 11073
rect 12110 11046 12194 11047
rect 12110 11041 12138 11046
rect 12166 10962 12194 11046
rect 12222 10962 12250 11942
rect 12278 11937 12306 11942
rect 12670 11914 12698 11919
rect 12334 11913 12698 11914
rect 12334 11887 12671 11913
rect 12697 11887 12698 11913
rect 12334 11886 12698 11887
rect 12278 11858 12306 11863
rect 12278 11633 12306 11830
rect 12278 11607 12279 11633
rect 12305 11607 12306 11633
rect 12278 11601 12306 11607
rect 12334 11521 12362 11886
rect 12670 11881 12698 11886
rect 12894 11914 12922 11919
rect 12334 11495 12335 11521
rect 12361 11495 12362 11521
rect 12334 11489 12362 11495
rect 12502 11690 12530 11695
rect 12278 10962 12306 10967
rect 12166 10934 12278 10962
rect 12278 10929 12306 10934
rect 12110 10906 12138 10911
rect 12110 10859 12138 10878
rect 11886 10457 12082 10458
rect 11886 10431 11887 10457
rect 11913 10431 12082 10457
rect 11886 10430 12082 10431
rect 12222 10793 12250 10799
rect 12222 10767 12223 10793
rect 12249 10767 12250 10793
rect 11774 10402 11802 10407
rect 11718 10374 11774 10402
rect 11774 10355 11802 10374
rect 11662 10094 11858 10122
rect 11494 9505 11522 9982
rect 11550 9618 11578 9623
rect 11774 9618 11802 9623
rect 11550 9617 11802 9618
rect 11550 9591 11551 9617
rect 11577 9591 11775 9617
rect 11801 9591 11802 9617
rect 11550 9590 11802 9591
rect 11550 9585 11578 9590
rect 11494 9479 11495 9505
rect 11521 9479 11522 9505
rect 11494 9473 11522 9479
rect 11438 9366 11522 9394
rect 11326 9338 11354 9343
rect 11326 9291 11354 9310
rect 11102 9226 11130 9231
rect 11102 9179 11130 9198
rect 11158 8834 11186 9254
rect 11438 9226 11466 9231
rect 11382 9198 11438 9226
rect 11270 9170 11298 9175
rect 11270 9123 11298 9142
rect 11382 8945 11410 9198
rect 11438 9179 11466 9198
rect 11438 9058 11466 9063
rect 11494 9058 11522 9366
rect 11606 9282 11634 9287
rect 11606 9235 11634 9254
rect 11466 9030 11522 9058
rect 11774 9225 11802 9590
rect 11774 9199 11775 9225
rect 11801 9199 11802 9225
rect 11438 9025 11466 9030
rect 11382 8919 11383 8945
rect 11409 8919 11410 8945
rect 11382 8913 11410 8919
rect 11774 8834 11802 9199
rect 11158 8833 11298 8834
rect 11158 8807 11159 8833
rect 11185 8807 11298 8833
rect 11158 8806 11298 8807
rect 11158 8801 11186 8806
rect 10766 8358 10934 8386
rect 10654 8050 10682 8055
rect 10654 8003 10682 8022
rect 10766 8049 10794 8358
rect 10934 8339 10962 8358
rect 11158 8721 11186 8727
rect 11158 8695 11159 8721
rect 11185 8695 11186 8721
rect 11158 8162 11186 8695
rect 11158 8129 11186 8134
rect 10766 8023 10767 8049
rect 10793 8023 10794 8049
rect 10318 7993 10374 7994
rect 10318 7967 10319 7993
rect 10345 7967 10374 7993
rect 10318 7966 10374 7967
rect 10318 7961 10346 7966
rect 10374 7947 10402 7966
rect 10430 7938 10458 7943
rect 10430 7891 10458 7910
rect 10710 7937 10738 7943
rect 10710 7911 10711 7937
rect 10737 7911 10738 7937
rect 10038 7769 10122 7770
rect 10038 7743 10039 7769
rect 10065 7743 10122 7769
rect 10038 7742 10122 7743
rect 10038 7737 10066 7742
rect 9758 7625 9786 7630
rect 9814 7713 9842 7719
rect 9814 7687 9815 7713
rect 9841 7687 9842 7713
rect 8806 7462 9002 7490
rect 8414 6903 8415 6929
rect 8441 6903 8442 6929
rect 8414 6897 8442 6903
rect 8918 7322 8946 7327
rect 8974 7322 9002 7462
rect 9030 7322 9058 7327
rect 8974 7321 9058 7322
rect 8974 7295 9031 7321
rect 9057 7295 9058 7321
rect 8974 7294 9058 7295
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 8918 6481 8946 7294
rect 8918 6455 8919 6481
rect 8945 6455 8946 6481
rect 8918 6449 8946 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 9030 4214 9058 7294
rect 9198 7322 9226 7574
rect 9814 7377 9842 7687
rect 10038 7658 10066 7663
rect 9982 7601 10010 7607
rect 9982 7575 9983 7601
rect 10009 7575 10010 7601
rect 9982 7574 10010 7575
rect 9814 7351 9815 7377
rect 9841 7351 9842 7377
rect 9814 7345 9842 7351
rect 9870 7546 10010 7574
rect 9254 7322 9282 7327
rect 9226 7321 9282 7322
rect 9226 7295 9255 7321
rect 9281 7295 9282 7321
rect 9226 7294 9282 7295
rect 9198 7275 9226 7294
rect 9254 7289 9282 7294
rect 9870 7266 9898 7546
rect 9310 7238 9898 7266
rect 9254 6538 9282 6543
rect 9310 6538 9338 7238
rect 10038 7210 10066 7630
rect 10710 7434 10738 7911
rect 10766 7770 10794 8023
rect 11270 8049 11298 8806
rect 11774 8801 11802 8806
rect 11438 8777 11466 8783
rect 11438 8751 11439 8777
rect 11465 8751 11466 8777
rect 11270 8023 11271 8049
rect 11297 8023 11298 8049
rect 11270 8017 11298 8023
rect 11382 8442 11410 8447
rect 11158 7994 11186 7999
rect 11158 7947 11186 7966
rect 10878 7938 10906 7943
rect 10878 7891 10906 7910
rect 10766 7737 10794 7742
rect 11382 7574 11410 8414
rect 9870 7182 10066 7210
rect 10486 7406 10738 7434
rect 11326 7546 11410 7574
rect 11438 8050 11466 8751
rect 11438 7574 11466 8022
rect 11606 8777 11634 8783
rect 11606 8751 11607 8777
rect 11633 8751 11634 8777
rect 11606 8106 11634 8751
rect 11494 7994 11522 7999
rect 11494 7947 11522 7966
rect 11606 7657 11634 8078
rect 11662 8386 11690 8391
rect 11830 8386 11858 10094
rect 11886 9898 11914 10430
rect 12222 9954 12250 10767
rect 12502 10738 12530 11662
rect 12782 11690 12810 11695
rect 12782 11643 12810 11662
rect 12838 11634 12866 11639
rect 12838 11587 12866 11606
rect 12614 11577 12642 11583
rect 12614 11551 12615 11577
rect 12641 11551 12642 11577
rect 12614 11354 12642 11551
rect 12614 11321 12642 11326
rect 12894 11577 12922 11886
rect 13734 11690 13762 11998
rect 13958 12025 13986 12670
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 13958 11999 13959 12025
rect 13985 11999 13986 12025
rect 13958 11993 13986 11999
rect 14070 12306 14098 12311
rect 14070 11969 14098 12278
rect 14462 12306 14490 12311
rect 14462 12259 14490 12278
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 14070 11943 14071 11969
rect 14097 11943 14098 11969
rect 14070 11937 14098 11943
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 13902 11914 13930 11919
rect 13902 11867 13930 11886
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 13734 11657 13762 11662
rect 12894 11551 12895 11577
rect 12921 11551 12922 11577
rect 12838 10962 12866 10967
rect 12726 10850 12754 10855
rect 12726 10793 12754 10822
rect 12726 10767 12727 10793
rect 12753 10767 12754 10793
rect 12726 10761 12754 10767
rect 12614 10738 12642 10743
rect 12502 10737 12642 10738
rect 12502 10711 12615 10737
rect 12641 10711 12642 10737
rect 12502 10710 12642 10711
rect 12278 10402 12306 10407
rect 12278 10355 12306 10374
rect 11886 9865 11914 9870
rect 12054 9926 12222 9954
rect 11998 9730 12026 9735
rect 11998 9683 12026 9702
rect 11886 9618 11914 9623
rect 11886 8833 11914 9590
rect 12054 9561 12082 9926
rect 12222 9921 12250 9926
rect 12502 9730 12530 10710
rect 12614 10705 12642 10710
rect 12502 9697 12530 9702
rect 12558 10458 12586 10463
rect 12558 10401 12586 10430
rect 12558 10375 12559 10401
rect 12585 10375 12586 10401
rect 12558 10066 12586 10375
rect 12838 10402 12866 10934
rect 12894 10906 12922 11551
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 12894 10873 12922 10878
rect 13622 10906 13650 10911
rect 13230 10849 13258 10855
rect 13230 10823 13231 10849
rect 13257 10823 13258 10849
rect 12894 10794 12922 10799
rect 13062 10794 13090 10799
rect 12894 10793 13090 10794
rect 12894 10767 12895 10793
rect 12921 10767 13063 10793
rect 13089 10767 13090 10793
rect 12894 10766 13090 10767
rect 12894 10761 12922 10766
rect 13062 10761 13090 10766
rect 13230 10457 13258 10823
rect 13230 10431 13231 10457
rect 13257 10431 13258 10457
rect 13230 10425 13258 10431
rect 12894 10402 12922 10407
rect 12838 10401 12922 10402
rect 12838 10375 12895 10401
rect 12921 10375 12922 10401
rect 12838 10374 12922 10375
rect 12894 10122 12922 10374
rect 12950 10122 12978 10127
rect 12894 10121 12978 10122
rect 12894 10095 12951 10121
rect 12977 10095 12978 10121
rect 12894 10094 12978 10095
rect 12950 10089 12978 10094
rect 12670 10066 12698 10071
rect 12558 10065 12698 10066
rect 12558 10039 12671 10065
rect 12697 10039 12698 10065
rect 12558 10038 12698 10039
rect 12222 9618 12250 9623
rect 12502 9618 12530 9623
rect 12558 9618 12586 10038
rect 12670 10033 12698 10038
rect 13118 10009 13146 10015
rect 13118 9983 13119 10009
rect 13145 9983 13146 10009
rect 12614 9954 12642 9959
rect 12614 9907 12642 9926
rect 12250 9590 12418 9618
rect 12222 9571 12250 9590
rect 12054 9535 12055 9561
rect 12081 9535 12082 9561
rect 12054 9338 12082 9535
rect 12054 9305 12082 9310
rect 11886 8807 11887 8833
rect 11913 8807 11914 8833
rect 11886 8801 11914 8807
rect 12054 8834 12082 8839
rect 12054 8787 12082 8806
rect 12390 8833 12418 9590
rect 12502 9617 12586 9618
rect 12502 9591 12503 9617
rect 12529 9591 12586 9617
rect 12502 9590 12586 9591
rect 12502 9585 12530 9590
rect 12782 9562 12810 9567
rect 12782 9337 12810 9534
rect 12782 9311 12783 9337
rect 12809 9311 12810 9337
rect 12782 9305 12810 9311
rect 12950 9506 12978 9511
rect 13118 9506 13146 9983
rect 13510 9954 13538 9959
rect 13454 9953 13538 9954
rect 13454 9927 13511 9953
rect 13537 9927 13538 9953
rect 13454 9926 13538 9927
rect 13230 9898 13258 9903
rect 13230 9617 13258 9870
rect 13230 9591 13231 9617
rect 13257 9591 13258 9617
rect 13230 9585 13258 9591
rect 13342 9562 13370 9567
rect 13342 9515 13370 9534
rect 12950 9505 13146 9506
rect 12950 9479 12951 9505
rect 12977 9479 13146 9505
rect 12950 9478 13146 9479
rect 13454 9505 13482 9926
rect 13510 9921 13538 9926
rect 13454 9479 13455 9505
rect 13481 9479 13482 9505
rect 12614 9226 12642 9231
rect 12614 9179 12642 9198
rect 12390 8807 12391 8833
rect 12417 8807 12418 8833
rect 12390 8801 12418 8807
rect 12726 8834 12754 8839
rect 12278 8722 12306 8727
rect 12278 8675 12306 8694
rect 11662 7993 11690 8358
rect 11662 7967 11663 7993
rect 11689 7967 11690 7993
rect 11662 7961 11690 7967
rect 11774 8358 11858 8386
rect 11774 8330 11802 8358
rect 11606 7631 11607 7657
rect 11633 7631 11634 7657
rect 11606 7625 11634 7631
rect 11774 7657 11802 8302
rect 12054 8162 12082 8167
rect 12054 8115 12082 8134
rect 12110 8106 12138 8111
rect 12110 8049 12138 8078
rect 12726 8105 12754 8806
rect 12782 8442 12810 8447
rect 12950 8442 12978 9478
rect 13454 9473 13482 9479
rect 13510 9729 13538 9735
rect 13510 9703 13511 9729
rect 13537 9703 13538 9729
rect 13510 9506 13538 9703
rect 13622 9617 13650 10878
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 14294 10458 14322 10463
rect 14294 10411 14322 10430
rect 18830 10010 18858 10015
rect 18830 9963 18858 9982
rect 13958 9954 13986 9959
rect 13846 9674 13874 9679
rect 13622 9591 13623 9617
rect 13649 9591 13650 9617
rect 13622 9585 13650 9591
rect 13678 9673 13874 9674
rect 13678 9647 13847 9673
rect 13873 9647 13874 9673
rect 13678 9646 13874 9647
rect 13678 9506 13706 9646
rect 13846 9641 13874 9646
rect 13958 9617 13986 9926
rect 14574 9954 14602 9959
rect 14574 9907 14602 9926
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 13958 9591 13959 9617
rect 13985 9591 13986 9617
rect 13958 9585 13986 9591
rect 13510 9478 13706 9506
rect 13790 9562 13818 9567
rect 12810 8441 12978 8442
rect 12810 8415 12951 8441
rect 12977 8415 12978 8441
rect 12810 8414 12978 8415
rect 12782 8395 12810 8414
rect 12726 8079 12727 8105
rect 12753 8079 12754 8105
rect 12726 8073 12754 8079
rect 12110 8023 12111 8049
rect 12137 8023 12138 8049
rect 12110 8017 12138 8023
rect 12502 8050 12530 8055
rect 12502 8003 12530 8022
rect 11830 7994 11858 7999
rect 11830 7947 11858 7966
rect 11942 7994 11970 7999
rect 11942 7947 11970 7966
rect 12726 7994 12754 7999
rect 11774 7631 11775 7657
rect 11801 7631 11802 7657
rect 11774 7625 11802 7631
rect 11886 7937 11914 7943
rect 11886 7911 11887 7937
rect 11913 7911 11914 7937
rect 11886 7657 11914 7911
rect 11886 7631 11887 7657
rect 11913 7631 11914 7657
rect 11886 7625 11914 7631
rect 11718 7601 11746 7607
rect 11718 7575 11719 7601
rect 11745 7575 11746 7601
rect 11718 7574 11746 7575
rect 11438 7546 11578 7574
rect 9870 7181 9898 7182
rect 9254 6537 9338 6538
rect 9254 6511 9255 6537
rect 9281 6511 9338 6537
rect 9254 6510 9338 6511
rect 9814 7153 9842 7159
rect 9814 7127 9815 7153
rect 9841 7127 9842 7153
rect 9870 7155 9871 7181
rect 9897 7155 9898 7181
rect 9870 7149 9898 7155
rect 9814 6538 9842 7127
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10486 6929 10514 7406
rect 10486 6903 10487 6929
rect 10513 6903 10514 6929
rect 10486 6897 10514 6903
rect 10766 7266 10794 7271
rect 10150 6874 10178 6879
rect 10150 6827 10178 6846
rect 10766 6874 10794 7238
rect 11326 7266 11354 7546
rect 11326 7219 11354 7238
rect 9254 6505 9282 6510
rect 9814 6505 9842 6510
rect 10318 6538 10346 6543
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 8806 4186 9058 4214
rect 10318 4214 10346 6510
rect 10766 6537 10794 6846
rect 11550 6817 11578 7546
rect 11662 7546 11746 7574
rect 11662 7321 11690 7546
rect 11662 7295 11663 7321
rect 11689 7295 11690 7321
rect 11662 7289 11690 7295
rect 12726 7321 12754 7966
rect 12894 7770 12922 8414
rect 12950 8409 12978 8414
rect 13230 8833 13258 8839
rect 13230 8807 13231 8833
rect 13257 8807 13258 8833
rect 13174 8162 13202 8167
rect 13230 8162 13258 8807
rect 13398 8777 13426 8783
rect 13398 8751 13399 8777
rect 13425 8751 13426 8777
rect 13202 8134 13258 8162
rect 13286 8722 13314 8727
rect 13174 8115 13202 8134
rect 12950 8106 12978 8111
rect 12950 8049 12978 8078
rect 12950 8023 12951 8049
rect 12977 8023 12978 8049
rect 12950 8017 12978 8023
rect 13062 8050 13090 8055
rect 13286 8050 13314 8694
rect 13342 8721 13370 8727
rect 13342 8695 13343 8721
rect 13369 8695 13370 8721
rect 13342 8497 13370 8695
rect 13342 8471 13343 8497
rect 13369 8471 13370 8497
rect 13342 8465 13370 8471
rect 13398 8330 13426 8751
rect 13398 8302 13650 8330
rect 13566 8218 13594 8223
rect 13342 8050 13370 8055
rect 13286 8049 13370 8050
rect 13286 8023 13343 8049
rect 13369 8023 13370 8049
rect 13286 8022 13370 8023
rect 13062 8003 13090 8022
rect 13342 8017 13370 8022
rect 13566 8049 13594 8190
rect 13622 8105 13650 8302
rect 13622 8079 13623 8105
rect 13649 8079 13650 8105
rect 13622 8073 13650 8079
rect 13566 8023 13567 8049
rect 13593 8023 13594 8049
rect 13566 8017 13594 8023
rect 13678 8050 13706 8055
rect 13790 8050 13818 9534
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 18942 8833 18970 8839
rect 18942 8807 18943 8833
rect 18969 8807 18970 8833
rect 18830 8442 18858 8447
rect 18774 8441 18858 8442
rect 18774 8415 18831 8441
rect 18857 8415 18858 8441
rect 18774 8414 18858 8415
rect 14406 8386 14434 8391
rect 14406 8218 14434 8358
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 14406 8185 14434 8190
rect 13846 8050 13874 8055
rect 13678 8049 13874 8050
rect 13678 8023 13679 8049
rect 13705 8023 13847 8049
rect 13873 8023 13874 8049
rect 13678 8022 13874 8023
rect 13678 8017 13706 8022
rect 13846 8017 13874 8022
rect 13902 8050 13930 8055
rect 13902 8003 13930 8022
rect 14014 8049 14042 8055
rect 14014 8023 14015 8049
rect 14041 8023 14042 8049
rect 13230 7994 13258 7999
rect 13230 7993 13314 7994
rect 13230 7967 13231 7993
rect 13257 7967 13314 7993
rect 13230 7966 13314 7967
rect 13230 7961 13258 7966
rect 12894 7769 13090 7770
rect 12894 7743 12895 7769
rect 12921 7743 13090 7769
rect 12894 7742 13090 7743
rect 12894 7737 12922 7742
rect 13062 7657 13090 7742
rect 13286 7714 13314 7966
rect 13454 7714 13482 7719
rect 13286 7713 13482 7714
rect 13286 7687 13455 7713
rect 13481 7687 13482 7713
rect 13286 7686 13482 7687
rect 13454 7681 13482 7686
rect 13062 7631 13063 7657
rect 13089 7631 13090 7657
rect 13062 7574 13090 7631
rect 14014 7658 14042 8023
rect 14854 7714 14882 7719
rect 14854 7667 14882 7686
rect 14742 7658 14770 7663
rect 14014 7625 14042 7630
rect 14518 7630 14742 7658
rect 14518 7601 14546 7630
rect 14518 7575 14519 7601
rect 14545 7575 14546 7601
rect 13062 7546 13314 7574
rect 14518 7569 14546 7575
rect 12726 7295 12727 7321
rect 12753 7295 12754 7321
rect 11774 7266 11802 7271
rect 11774 6985 11802 7238
rect 11774 6959 11775 6985
rect 11801 6959 11802 6985
rect 11774 6953 11802 6959
rect 12726 7154 12754 7295
rect 13286 7321 13314 7546
rect 13286 7295 13287 7321
rect 13313 7295 13314 7321
rect 13286 7289 13314 7295
rect 14630 7265 14658 7630
rect 14742 7611 14770 7630
rect 18774 7658 18802 8414
rect 18830 8409 18858 8414
rect 18942 8386 18970 8807
rect 20006 8442 20034 8863
rect 20006 8409 20034 8414
rect 18942 8353 18970 8358
rect 19950 8385 19978 8391
rect 19950 8359 19951 8385
rect 19977 8359 19978 8385
rect 19950 8106 19978 8359
rect 19950 8073 19978 8078
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 18830 7770 18858 8023
rect 18830 7737 18858 7742
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18774 7625 18802 7630
rect 18830 7657 18858 7663
rect 18830 7631 18831 7657
rect 18857 7631 18858 7657
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 14630 7239 14631 7265
rect 14657 7239 14658 7265
rect 14630 7233 14658 7239
rect 12894 7154 12922 7159
rect 12726 7153 12922 7154
rect 12726 7127 12895 7153
rect 12921 7127 12922 7153
rect 12726 7126 12922 7127
rect 11550 6791 11551 6817
rect 11577 6791 11578 6817
rect 11550 6785 11578 6791
rect 10766 6511 10767 6537
rect 10793 6511 10794 6537
rect 10766 6505 10794 6511
rect 12726 4214 12754 7126
rect 12894 7121 12922 7126
rect 13062 7153 13090 7159
rect 13062 7127 13063 7153
rect 13089 7127 13090 7153
rect 13062 4214 13090 7127
rect 14742 7154 14770 7159
rect 14742 7107 14770 7126
rect 18830 7154 18858 7631
rect 20006 7601 20034 7607
rect 20006 7575 20007 7601
rect 20033 7575 20034 7601
rect 20006 7434 20034 7575
rect 20006 7401 20034 7406
rect 18830 7121 18858 7126
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 10318 4186 10402 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8806 1777 8834 4186
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 10374 1777 10402 4186
rect 12614 4186 12754 4214
rect 12894 4186 13090 4214
rect 10374 1751 10375 1777
rect 10401 1751 10402 1777
rect 10374 1745 10402 1751
rect 12446 1834 12474 1839
rect 10094 1722 10122 1727
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10094 400 10122 1694
rect 10878 1722 10906 1727
rect 10878 1665 10906 1694
rect 12278 1666 12306 1671
rect 10878 1639 10879 1665
rect 10905 1639 10906 1665
rect 10878 1633 10906 1639
rect 12110 1665 12306 1666
rect 12110 1639 12279 1665
rect 12305 1639 12306 1665
rect 12110 1638 12306 1639
rect 12110 400 12138 1638
rect 12278 1633 12306 1638
rect 12446 400 12474 1806
rect 12614 1777 12642 4186
rect 12894 2169 12922 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12894 2143 12895 2169
rect 12921 2143 12922 2169
rect 12894 2137 12922 2143
rect 12614 1751 12615 1777
rect 12641 1751 12642 1777
rect 12614 1745 12642 1751
rect 12782 2058 12810 2063
rect 12782 400 12810 2030
rect 13398 2058 13426 2063
rect 13398 2011 13426 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 13062 1834 13090 1839
rect 13062 1787 13090 1806
rect 9072 0 9128 400
rect 10080 0 10136 400
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 12782 19278 12810 19306
rect 13398 19278 13426 19306
rect 11774 19110 11802 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 10094 18718 10122 18746
rect 10710 18745 10738 18746
rect 10710 18719 10711 18745
rect 10711 18719 10737 18745
rect 10737 18719 10738 18745
rect 10710 18718 10738 18719
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 2086 13790 2114 13818
rect 966 13118 994 13146
rect 966 12782 994 12810
rect 966 11774 994 11802
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 966 10737 994 10738
rect 966 10711 967 10737
rect 967 10711 993 10737
rect 993 10711 994 10737
rect 966 10710 994 10711
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2142 13537 2170 13538
rect 2142 13511 2143 13537
rect 2143 13511 2169 13537
rect 2169 13511 2170 13537
rect 2142 13510 2170 13511
rect 6174 13510 6202 13538
rect 7126 13230 7154 13258
rect 6174 13174 6202 13202
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 6062 13118 6090 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 7126 12670 7154 12698
rect 7350 12894 7378 12922
rect 7798 13398 7826 13426
rect 7630 13257 7658 13258
rect 7630 13231 7631 13257
rect 7631 13231 7657 13257
rect 7657 13231 7658 13257
rect 7630 13230 7658 13231
rect 7742 13201 7770 13202
rect 7742 13175 7743 13201
rect 7743 13175 7769 13201
rect 7769 13175 7770 13201
rect 7742 13174 7770 13175
rect 7574 13118 7602 13146
rect 8190 13118 8218 13146
rect 8694 13145 8722 13146
rect 8694 13119 8695 13145
rect 8695 13119 8721 13145
rect 8721 13119 8722 13145
rect 8694 13118 8722 13119
rect 7462 12697 7490 12698
rect 7462 12671 7463 12697
rect 7463 12671 7489 12697
rect 7489 12671 7490 12697
rect 7462 12670 7490 12671
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 6902 11969 6930 11970
rect 6902 11943 6903 11969
rect 6903 11943 6929 11969
rect 6929 11943 6930 11969
rect 6902 11942 6930 11943
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 5334 11521 5362 11522
rect 5334 11495 5335 11521
rect 5335 11495 5361 11521
rect 5361 11495 5362 11521
rect 5334 11494 5362 11495
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 6398 11102 6426 11130
rect 6622 11158 6650 11186
rect 5334 10990 5362 11018
rect 2142 10793 2170 10794
rect 2142 10767 2143 10793
rect 2143 10767 2169 10793
rect 2169 10767 2170 10793
rect 2142 10766 2170 10767
rect 5222 10766 5250 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6286 10737 6314 10738
rect 6286 10711 6287 10737
rect 6287 10711 6313 10737
rect 6313 10711 6314 10737
rect 6286 10710 6314 10711
rect 6734 11129 6762 11130
rect 6734 11103 6735 11129
rect 6735 11103 6761 11129
rect 6761 11103 6762 11129
rect 6734 11102 6762 11103
rect 6958 11886 6986 11914
rect 6958 11521 6986 11522
rect 6958 11495 6959 11521
rect 6959 11495 6985 11521
rect 6985 11495 6986 11521
rect 6958 11494 6986 11495
rect 7406 11438 7434 11466
rect 7462 12558 7490 12586
rect 6958 11382 6986 11410
rect 6902 11129 6930 11130
rect 6902 11103 6903 11129
rect 6903 11103 6929 11129
rect 6929 11103 6930 11129
rect 6902 11102 6930 11103
rect 6790 10878 6818 10906
rect 7126 10878 7154 10906
rect 5222 10374 5250 10402
rect 2086 10262 2114 10290
rect 6902 10737 6930 10738
rect 6902 10711 6903 10737
rect 6903 10711 6929 10737
rect 6929 10711 6930 10737
rect 6902 10710 6930 10711
rect 6902 10401 6930 10402
rect 6902 10375 6903 10401
rect 6903 10375 6929 10401
rect 6929 10375 6930 10401
rect 6902 10374 6930 10375
rect 7686 12753 7714 12754
rect 7686 12727 7687 12753
rect 7687 12727 7713 12753
rect 7713 12727 7714 12753
rect 7686 12726 7714 12727
rect 7630 12278 7658 12306
rect 7854 12305 7882 12306
rect 7854 12279 7855 12305
rect 7855 12279 7881 12305
rect 7881 12279 7882 12305
rect 7854 12278 7882 12279
rect 8694 12278 8722 12306
rect 7630 11942 7658 11970
rect 7910 11886 7938 11914
rect 7574 11270 7602 11298
rect 7686 11438 7714 11466
rect 8358 11886 8386 11914
rect 8022 11830 8050 11858
rect 8470 11857 8498 11858
rect 8470 11831 8471 11857
rect 8471 11831 8497 11857
rect 8497 11831 8498 11857
rect 8470 11830 8498 11831
rect 8918 12278 8946 12306
rect 8582 11606 8610 11634
rect 8694 11718 8722 11746
rect 8582 11494 8610 11522
rect 7966 11297 7994 11298
rect 7966 11271 7967 11297
rect 7967 11271 7993 11297
rect 7993 11271 7994 11297
rect 7966 11270 7994 11271
rect 7630 11129 7658 11130
rect 7630 11103 7631 11129
rect 7631 11103 7657 11129
rect 7657 11103 7658 11129
rect 7630 11102 7658 11103
rect 7630 10990 7658 11018
rect 8694 11382 8722 11410
rect 9030 13929 9058 13930
rect 9030 13903 9031 13929
rect 9031 13903 9057 13929
rect 9057 13903 9058 13929
rect 9030 13902 9058 13903
rect 9366 13929 9394 13930
rect 9366 13903 9367 13929
rect 9367 13903 9393 13929
rect 9393 13903 9394 13929
rect 9366 13902 9394 13903
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9870 13929 9898 13930
rect 9870 13903 9871 13929
rect 9871 13903 9897 13929
rect 9897 13903 9898 13929
rect 9870 13902 9898 13903
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 10822 13846 10850 13874
rect 9870 13510 9898 13538
rect 9534 13230 9562 13258
rect 10206 13510 10234 13538
rect 9086 12726 9114 12754
rect 8974 11550 9002 11578
rect 8862 11465 8890 11466
rect 8862 11439 8863 11465
rect 8863 11439 8889 11465
rect 8889 11439 8890 11465
rect 8862 11438 8890 11439
rect 8806 11185 8834 11186
rect 8806 11159 8807 11185
rect 8807 11159 8833 11185
rect 8833 11159 8834 11185
rect 8806 11158 8834 11159
rect 9030 11606 9058 11634
rect 8806 11046 8834 11074
rect 7350 10374 7378 10402
rect 6342 10065 6370 10066
rect 6342 10039 6343 10065
rect 6343 10039 6369 10065
rect 6369 10039 6370 10065
rect 6342 10038 6370 10039
rect 6846 10038 6874 10066
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 7406 9982 7434 10010
rect 6902 9870 6930 9898
rect 7294 9478 7322 9506
rect 6006 9198 6034 9226
rect 6398 9142 6426 9170
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 5614 8806 5642 8834
rect 966 8078 994 8106
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 7126 9169 7154 9170
rect 7126 9143 7127 9169
rect 7127 9143 7153 9169
rect 7153 9143 7154 9169
rect 7126 9142 7154 9143
rect 7182 8806 7210 8834
rect 7966 10793 7994 10794
rect 7966 10767 7967 10793
rect 7967 10767 7993 10793
rect 7993 10767 7994 10793
rect 7966 10766 7994 10767
rect 7854 10094 7882 10122
rect 8022 10430 8050 10458
rect 8638 10457 8666 10458
rect 8638 10431 8639 10457
rect 8639 10431 8665 10457
rect 8665 10431 8666 10457
rect 8638 10430 8666 10431
rect 8526 10094 8554 10122
rect 9030 11158 9058 11186
rect 8974 11102 9002 11130
rect 8750 10793 8778 10794
rect 8750 10767 8751 10793
rect 8751 10767 8777 10793
rect 8777 10767 8778 10793
rect 8750 10766 8778 10767
rect 7966 9897 7994 9898
rect 7966 9871 7967 9897
rect 7967 9871 7993 9897
rect 7993 9871 7994 9897
rect 7966 9870 7994 9871
rect 8134 9897 8162 9898
rect 8134 9871 8135 9897
rect 8135 9871 8161 9897
rect 8161 9871 8162 9897
rect 8134 9870 8162 9871
rect 7742 9478 7770 9506
rect 8470 10038 8498 10066
rect 8414 9926 8442 9954
rect 8358 9870 8386 9898
rect 8246 9478 8274 9506
rect 8694 10009 8722 10010
rect 8694 9983 8695 10009
rect 8695 9983 8721 10009
rect 8721 9983 8722 10009
rect 8694 9982 8722 9983
rect 8750 9814 8778 9842
rect 8862 9814 8890 9842
rect 7518 9198 7546 9226
rect 7350 9030 7378 9058
rect 7014 8358 7042 8386
rect 7574 8358 7602 8386
rect 2142 7574 2170 7602
rect 5894 7601 5922 7602
rect 5894 7575 5895 7601
rect 5895 7575 5921 7601
rect 5921 7575 5922 7601
rect 5894 7574 5922 7575
rect 7014 7910 7042 7938
rect 7910 8694 7938 8722
rect 8358 8721 8386 8722
rect 8358 8695 8359 8721
rect 8359 8695 8385 8721
rect 8385 8695 8386 8721
rect 8358 8694 8386 8695
rect 8582 9310 8610 9338
rect 8918 9478 8946 9506
rect 9254 12726 9282 12754
rect 9814 13398 9842 13426
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9814 12753 9842 12754
rect 9814 12727 9815 12753
rect 9815 12727 9841 12753
rect 9841 12727 9842 12753
rect 9814 12726 9842 12727
rect 9926 13230 9954 13258
rect 11326 13873 11354 13874
rect 11326 13847 11327 13873
rect 11327 13847 11353 13873
rect 11353 13847 11354 13873
rect 11326 13846 11354 13847
rect 10878 13481 10906 13482
rect 10878 13455 10879 13481
rect 10879 13455 10905 13481
rect 10905 13455 10906 13481
rect 10878 13454 10906 13455
rect 9310 11577 9338 11578
rect 9310 11551 9311 11577
rect 9311 11551 9337 11577
rect 9337 11551 9338 11577
rect 9310 11550 9338 11551
rect 9198 11326 9226 11354
rect 9086 11073 9114 11074
rect 9086 11047 9087 11073
rect 9087 11047 9113 11073
rect 9113 11047 9114 11073
rect 9086 11046 9114 11047
rect 9198 10822 9226 10850
rect 9142 10766 9170 10794
rect 9086 10401 9114 10402
rect 9086 10375 9087 10401
rect 9087 10375 9113 10401
rect 9113 10375 9114 10401
rect 9086 10374 9114 10375
rect 9030 9982 9058 10010
rect 9198 10065 9226 10066
rect 9198 10039 9199 10065
rect 9199 10039 9225 10065
rect 9225 10039 9226 10065
rect 9198 10038 9226 10039
rect 9142 9982 9170 10010
rect 8974 9310 9002 9338
rect 9030 9198 9058 9226
rect 8862 8638 8890 8666
rect 9254 9534 9282 9562
rect 9310 9478 9338 9506
rect 9590 11662 9618 11690
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9646 11606 9674 11634
rect 9758 11270 9786 11298
rect 9702 10793 9730 10794
rect 9702 10767 9703 10793
rect 9703 10767 9729 10793
rect 9729 10767 9730 10793
rect 9702 10766 9730 10767
rect 9646 10430 9674 10458
rect 9478 10289 9506 10290
rect 9478 10263 9479 10289
rect 9479 10263 9505 10289
rect 9505 10263 9506 10289
rect 9478 10262 9506 10263
rect 9422 10038 9450 10066
rect 9478 9897 9506 9898
rect 9478 9871 9479 9897
rect 9479 9871 9505 9897
rect 9505 9871 9506 9897
rect 9478 9870 9506 9871
rect 9142 9225 9170 9226
rect 9142 9199 9143 9225
rect 9143 9199 9169 9225
rect 9169 9199 9170 9225
rect 9142 9198 9170 9199
rect 9366 9198 9394 9226
rect 9534 9198 9562 9226
rect 9646 10262 9674 10290
rect 9926 11913 9954 11914
rect 9926 11887 9927 11913
rect 9927 11887 9953 11913
rect 9953 11887 9954 11913
rect 9926 11886 9954 11887
rect 9870 11830 9898 11858
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10374 13286 10402 13314
rect 11998 13398 12026 13426
rect 10374 12278 10402 12306
rect 10710 12278 10738 12306
rect 11494 12278 11522 12306
rect 11550 13118 11578 13146
rect 11550 12614 11578 12642
rect 10318 11662 10346 11690
rect 10990 11886 11018 11914
rect 10206 11577 10234 11578
rect 10206 11551 10207 11577
rect 10207 11551 10233 11577
rect 10233 11551 10234 11577
rect 10206 11550 10234 11551
rect 10038 11521 10066 11522
rect 10038 11495 10039 11521
rect 10039 11495 10065 11521
rect 10065 11495 10066 11521
rect 10038 11494 10066 11495
rect 10150 11241 10178 11242
rect 10150 11215 10151 11241
rect 10151 11215 10177 11241
rect 10177 11215 10178 11241
rect 10150 11214 10178 11215
rect 10262 11521 10290 11522
rect 10262 11495 10263 11521
rect 10263 11495 10289 11521
rect 10289 11495 10290 11521
rect 10262 11494 10290 11495
rect 10318 11382 10346 11410
rect 10262 11185 10290 11186
rect 10262 11159 10263 11185
rect 10263 11159 10289 11185
rect 10289 11159 10290 11185
rect 10262 11158 10290 11159
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9870 10766 9898 10794
rect 9870 10401 9898 10402
rect 9870 10375 9871 10401
rect 9871 10375 9897 10401
rect 9897 10375 9898 10401
rect 9870 10374 9898 10375
rect 10374 10849 10402 10850
rect 10374 10823 10375 10849
rect 10375 10823 10401 10849
rect 10401 10823 10402 10849
rect 10374 10822 10402 10823
rect 10318 10374 10346 10402
rect 10598 11577 10626 11578
rect 10598 11551 10599 11577
rect 10599 11551 10625 11577
rect 10625 11551 10626 11577
rect 10598 11550 10626 11551
rect 10710 11326 10738 11354
rect 10654 11214 10682 11242
rect 10542 10878 10570 10906
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9814 10038 9842 10066
rect 9646 9505 9674 9506
rect 9646 9479 9647 9505
rect 9647 9479 9673 9505
rect 9673 9479 9674 9505
rect 9646 9478 9674 9479
rect 9646 9254 9674 9282
rect 9590 8806 9618 8834
rect 9310 8694 9338 8722
rect 9534 8694 9562 8722
rect 8750 8302 8778 8330
rect 8918 8414 8946 8442
rect 6846 7574 6874 7602
rect 7574 7574 7602 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 10262 9814 10290 9842
rect 10206 9729 10234 9730
rect 10206 9703 10207 9729
rect 10207 9703 10233 9729
rect 10233 9703 10234 9729
rect 10206 9702 10234 9703
rect 10150 9534 10178 9562
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9814 9310 9842 9338
rect 10598 9758 10626 9786
rect 11046 11550 11074 11578
rect 10878 11465 10906 11466
rect 10878 11439 10879 11465
rect 10879 11439 10905 11465
rect 10905 11439 10906 11465
rect 10878 11438 10906 11439
rect 10934 10542 10962 10570
rect 10990 10401 11018 10402
rect 10990 10375 10991 10401
rect 10991 10375 11017 10401
rect 11017 10375 11018 10401
rect 10990 10374 11018 10375
rect 10934 10065 10962 10066
rect 10934 10039 10935 10065
rect 10935 10039 10961 10065
rect 10961 10039 10962 10065
rect 10934 10038 10962 10039
rect 10878 9702 10906 9730
rect 9030 8302 9058 8330
rect 8750 7657 8778 7658
rect 8750 7631 8751 7657
rect 8751 7631 8777 7657
rect 8777 7631 8778 7657
rect 8750 7630 8778 7631
rect 10094 9281 10122 9282
rect 10094 9255 10095 9281
rect 10095 9255 10121 9281
rect 10121 9255 10122 9281
rect 10094 9254 10122 9255
rect 9870 9225 9898 9226
rect 9870 9199 9871 9225
rect 9871 9199 9897 9225
rect 9897 9199 9898 9225
rect 9870 9198 9898 9199
rect 9814 8833 9842 8834
rect 9814 8807 9815 8833
rect 9815 8807 9841 8833
rect 9841 8807 9842 8833
rect 9814 8806 9842 8807
rect 9870 8721 9898 8722
rect 9870 8695 9871 8721
rect 9871 8695 9897 8721
rect 9897 8695 9898 8721
rect 9870 8694 9898 8695
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10150 8721 10178 8722
rect 10150 8695 10151 8721
rect 10151 8695 10177 8721
rect 10177 8695 10178 8721
rect 10150 8694 10178 8695
rect 10094 8022 10122 8050
rect 10822 9310 10850 9338
rect 10654 9254 10682 9282
rect 11102 11382 11130 11410
rect 11158 11494 11186 11522
rect 11606 11718 11634 11746
rect 11494 11438 11522 11466
rect 11774 13145 11802 13146
rect 11774 13119 11775 13145
rect 11775 13119 11801 13145
rect 11801 13119 11802 13145
rect 11774 13118 11802 13119
rect 11886 13145 11914 13146
rect 11886 13119 11887 13145
rect 11887 13119 11913 13145
rect 11913 13119 11914 13145
rect 11886 13118 11914 13119
rect 11998 11830 12026 11858
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12614 13145 12642 13146
rect 12614 13119 12615 13145
rect 12615 13119 12641 13145
rect 12641 13119 12642 13145
rect 12614 13118 12642 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 13286 12614 13314 12642
rect 12166 12278 12194 12306
rect 12670 12305 12698 12306
rect 12670 12279 12671 12305
rect 12671 12279 12697 12305
rect 12697 12279 12698 12305
rect 12670 12278 12698 12279
rect 13006 12278 13034 12306
rect 13734 12025 13762 12026
rect 13734 11999 13735 12025
rect 13735 11999 13761 12025
rect 13761 11999 13762 12025
rect 13734 11998 13762 11999
rect 12054 11718 12082 11746
rect 11830 11606 11858 11634
rect 12054 11633 12082 11634
rect 12054 11607 12055 11633
rect 12055 11607 12081 11633
rect 12081 11607 12082 11633
rect 12054 11606 12082 11607
rect 11214 10710 11242 10738
rect 11214 10457 11242 10458
rect 11214 10431 11215 10457
rect 11215 10431 11241 10457
rect 11241 10431 11242 10457
rect 11214 10430 11242 10431
rect 11102 9758 11130 9786
rect 10262 8777 10290 8778
rect 10262 8751 10263 8777
rect 10263 8751 10289 8777
rect 10289 8751 10290 8777
rect 10262 8750 10290 8751
rect 10710 8777 10738 8778
rect 10710 8751 10711 8777
rect 10711 8751 10737 8777
rect 10737 8751 10738 8777
rect 10710 8750 10738 8751
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9926 7769 9954 7770
rect 9926 7743 9927 7769
rect 9927 7743 9953 7769
rect 9953 7743 9954 7769
rect 9926 7742 9954 7743
rect 11494 10737 11522 10738
rect 11494 10711 11495 10737
rect 11495 10711 11521 10737
rect 11521 10711 11522 10737
rect 11494 10710 11522 10711
rect 11942 10849 11970 10850
rect 11942 10823 11943 10849
rect 11943 10823 11969 10849
rect 11969 10823 11970 10849
rect 11942 10822 11970 10823
rect 11326 9617 11354 9618
rect 11326 9591 11327 9617
rect 11327 9591 11353 9617
rect 11353 9591 11354 9617
rect 11326 9590 11354 9591
rect 11606 10542 11634 10570
rect 12278 11830 12306 11858
rect 12894 11886 12922 11914
rect 12502 11662 12530 11690
rect 12278 10934 12306 10962
rect 12110 10905 12138 10906
rect 12110 10879 12111 10905
rect 12111 10879 12137 10905
rect 12137 10879 12138 10905
rect 12110 10878 12138 10879
rect 11774 10401 11802 10402
rect 11774 10375 11775 10401
rect 11775 10375 11801 10401
rect 11801 10375 11802 10401
rect 11774 10374 11802 10375
rect 11494 9982 11522 10010
rect 11326 9337 11354 9338
rect 11326 9311 11327 9337
rect 11327 9311 11353 9337
rect 11353 9311 11354 9337
rect 11326 9310 11354 9311
rect 11158 9254 11186 9282
rect 11102 9225 11130 9226
rect 11102 9199 11103 9225
rect 11103 9199 11129 9225
rect 11129 9199 11130 9225
rect 11102 9198 11130 9199
rect 11438 9225 11466 9226
rect 11438 9199 11439 9225
rect 11439 9199 11465 9225
rect 11465 9199 11466 9225
rect 11438 9198 11466 9199
rect 11270 9169 11298 9170
rect 11270 9143 11271 9169
rect 11271 9143 11297 9169
rect 11297 9143 11298 9169
rect 11270 9142 11298 9143
rect 11606 9281 11634 9282
rect 11606 9255 11607 9281
rect 11607 9255 11633 9281
rect 11633 9255 11634 9281
rect 11606 9254 11634 9255
rect 11438 9030 11466 9058
rect 10934 8358 10962 8386
rect 10654 8049 10682 8050
rect 10654 8023 10655 8049
rect 10655 8023 10681 8049
rect 10681 8023 10682 8049
rect 10654 8022 10682 8023
rect 11158 8134 11186 8162
rect 10374 7966 10402 7994
rect 10430 7937 10458 7938
rect 10430 7911 10431 7937
rect 10431 7911 10457 7937
rect 10457 7911 10458 7937
rect 10430 7910 10458 7911
rect 9758 7630 9786 7658
rect 9198 7574 9226 7602
rect 8918 7294 8946 7322
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 10038 7630 10066 7658
rect 9198 7294 9226 7322
rect 11774 8806 11802 8834
rect 11382 8441 11410 8442
rect 11382 8415 11383 8441
rect 11383 8415 11409 8441
rect 11409 8415 11410 8441
rect 11382 8414 11410 8415
rect 11158 7993 11186 7994
rect 11158 7967 11159 7993
rect 11159 7967 11185 7993
rect 11185 7967 11186 7993
rect 11158 7966 11186 7967
rect 10878 7937 10906 7938
rect 10878 7911 10879 7937
rect 10879 7911 10905 7937
rect 10905 7911 10906 7937
rect 10878 7910 10906 7911
rect 10766 7742 10794 7770
rect 11438 8022 11466 8050
rect 11606 8078 11634 8106
rect 11494 7993 11522 7994
rect 11494 7967 11495 7993
rect 11495 7967 11521 7993
rect 11521 7967 11522 7993
rect 11494 7966 11522 7967
rect 12782 11689 12810 11690
rect 12782 11663 12783 11689
rect 12783 11663 12809 11689
rect 12809 11663 12810 11689
rect 12782 11662 12810 11663
rect 12838 11633 12866 11634
rect 12838 11607 12839 11633
rect 12839 11607 12865 11633
rect 12865 11607 12866 11633
rect 12838 11606 12866 11607
rect 12614 11326 12642 11354
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 14070 12278 14098 12306
rect 14462 12305 14490 12306
rect 14462 12279 14463 12305
rect 14463 12279 14489 12305
rect 14489 12279 14490 12305
rect 14462 12278 14490 12279
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 13902 11913 13930 11914
rect 13902 11887 13903 11913
rect 13903 11887 13929 11913
rect 13929 11887 13930 11913
rect 13902 11886 13930 11887
rect 20006 11774 20034 11802
rect 13734 11662 13762 11690
rect 12838 10934 12866 10962
rect 12726 10822 12754 10850
rect 12278 10401 12306 10402
rect 12278 10375 12279 10401
rect 12279 10375 12305 10401
rect 12305 10375 12306 10401
rect 12278 10374 12306 10375
rect 11886 9870 11914 9898
rect 12222 9926 12250 9954
rect 11998 9729 12026 9730
rect 11998 9703 11999 9729
rect 11999 9703 12025 9729
rect 12025 9703 12026 9729
rect 11998 9702 12026 9703
rect 11886 9590 11914 9618
rect 12502 9702 12530 9730
rect 12558 10430 12586 10458
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 12894 10878 12922 10906
rect 13622 10878 13650 10906
rect 12614 9953 12642 9954
rect 12614 9927 12615 9953
rect 12615 9927 12641 9953
rect 12641 9927 12642 9953
rect 12614 9926 12642 9927
rect 12222 9617 12250 9618
rect 12222 9591 12223 9617
rect 12223 9591 12249 9617
rect 12249 9591 12250 9617
rect 12222 9590 12250 9591
rect 12054 9310 12082 9338
rect 12054 8833 12082 8834
rect 12054 8807 12055 8833
rect 12055 8807 12081 8833
rect 12081 8807 12082 8833
rect 12054 8806 12082 8807
rect 12782 9534 12810 9562
rect 13230 9870 13258 9898
rect 13342 9561 13370 9562
rect 13342 9535 13343 9561
rect 13343 9535 13369 9561
rect 13369 9535 13370 9561
rect 13342 9534 13370 9535
rect 12614 9225 12642 9226
rect 12614 9199 12615 9225
rect 12615 9199 12641 9225
rect 12641 9199 12642 9225
rect 12614 9198 12642 9199
rect 12726 8806 12754 8834
rect 12278 8721 12306 8722
rect 12278 8695 12279 8721
rect 12279 8695 12305 8721
rect 12305 8695 12306 8721
rect 12278 8694 12306 8695
rect 11662 8358 11690 8386
rect 11774 8302 11802 8330
rect 12054 8161 12082 8162
rect 12054 8135 12055 8161
rect 12055 8135 12081 8161
rect 12081 8135 12082 8161
rect 12054 8134 12082 8135
rect 12110 8078 12138 8106
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 14294 10457 14322 10458
rect 14294 10431 14295 10457
rect 14295 10431 14321 10457
rect 14321 10431 14322 10457
rect 14294 10430 14322 10431
rect 18830 10009 18858 10010
rect 18830 9983 18831 10009
rect 18831 9983 18857 10009
rect 18857 9983 18858 10009
rect 18830 9982 18858 9983
rect 13958 9926 13986 9954
rect 14574 9953 14602 9954
rect 14574 9927 14575 9953
rect 14575 9927 14601 9953
rect 14601 9927 14602 9953
rect 14574 9926 14602 9927
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 9758 20034 9786
rect 13790 9561 13818 9562
rect 13790 9535 13791 9561
rect 13791 9535 13817 9561
rect 13817 9535 13818 9561
rect 13790 9534 13818 9535
rect 12782 8441 12810 8442
rect 12782 8415 12783 8441
rect 12783 8415 12809 8441
rect 12809 8415 12810 8441
rect 12782 8414 12810 8415
rect 12502 8049 12530 8050
rect 12502 8023 12503 8049
rect 12503 8023 12529 8049
rect 12529 8023 12530 8049
rect 12502 8022 12530 8023
rect 11830 7993 11858 7994
rect 11830 7967 11831 7993
rect 11831 7967 11857 7993
rect 11857 7967 11858 7993
rect 11830 7966 11858 7967
rect 11942 7993 11970 7994
rect 11942 7967 11943 7993
rect 11943 7967 11969 7993
rect 11969 7967 11970 7993
rect 11942 7966 11970 7967
rect 12726 7966 12754 7994
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10766 7238 10794 7266
rect 10150 6873 10178 6874
rect 10150 6847 10151 6873
rect 10151 6847 10177 6873
rect 10177 6847 10178 6873
rect 10150 6846 10178 6847
rect 11326 7265 11354 7266
rect 11326 7239 11327 7265
rect 11327 7239 11353 7265
rect 11353 7239 11354 7265
rect 11326 7238 11354 7239
rect 10766 6846 10794 6874
rect 9814 6510 9842 6538
rect 10318 6537 10346 6538
rect 10318 6511 10319 6537
rect 10319 6511 10345 6537
rect 10345 6511 10346 6537
rect 10318 6510 10346 6511
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 13174 8161 13202 8162
rect 13174 8135 13175 8161
rect 13175 8135 13201 8161
rect 13201 8135 13202 8161
rect 13174 8134 13202 8135
rect 13286 8694 13314 8722
rect 12950 8078 12978 8106
rect 13062 8049 13090 8050
rect 13062 8023 13063 8049
rect 13063 8023 13089 8049
rect 13089 8023 13090 8049
rect 13062 8022 13090 8023
rect 13566 8190 13594 8218
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14406 8385 14434 8386
rect 14406 8359 14407 8385
rect 14407 8359 14433 8385
rect 14433 8359 14434 8385
rect 14406 8358 14434 8359
rect 14406 8190 14434 8218
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 13902 8049 13930 8050
rect 13902 8023 13903 8049
rect 13903 8023 13929 8049
rect 13929 8023 13930 8049
rect 13902 8022 13930 8023
rect 14854 7713 14882 7714
rect 14854 7687 14855 7713
rect 14855 7687 14881 7713
rect 14881 7687 14882 7713
rect 14854 7686 14882 7687
rect 14014 7630 14042 7658
rect 14742 7657 14770 7658
rect 14742 7631 14743 7657
rect 14743 7631 14769 7657
rect 14769 7631 14770 7657
rect 14742 7630 14770 7631
rect 11774 7238 11802 7266
rect 20006 8414 20034 8442
rect 18942 8358 18970 8386
rect 19950 8078 19978 8106
rect 18830 7742 18858 7770
rect 20006 7742 20034 7770
rect 18774 7630 18802 7658
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 14742 7153 14770 7154
rect 14742 7127 14743 7153
rect 14743 7127 14769 7153
rect 14769 7127 14770 7153
rect 14742 7126 14770 7127
rect 20006 7406 20034 7434
rect 18830 7126 18858 7154
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 12446 1806 12474 1834
rect 10094 1694 10122 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 10878 1694 10906 1722
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12782 2030 12810 2058
rect 13398 2057 13426 2058
rect 13398 2031 13399 2057
rect 13399 2031 13425 2057
rect 13425 2031 13426 2057
rect 13398 2030 13426 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 13062 1833 13090 1834
rect 13062 1807 13063 1833
rect 13063 1807 13089 1833
rect 13089 1807 13090 1833
rect 13062 1806 13090 1807
<< metal3 >>
rect 12777 19278 12782 19306
rect 12810 19278 13398 19306
rect 13426 19278 13431 19306
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10089 18718 10094 18746
rect 10122 18718 10710 18746
rect 10738 18718 10743 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 9025 13902 9030 13930
rect 9058 13902 9366 13930
rect 9394 13902 9399 13930
rect 9865 13902 9870 13930
rect 9898 13902 10402 13930
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 2137 13510 2142 13538
rect 2170 13510 6174 13538
rect 6202 13510 6207 13538
rect 9865 13510 9870 13538
rect 9898 13510 10206 13538
rect 10234 13510 10239 13538
rect 7793 13398 7798 13426
rect 7826 13398 9814 13426
rect 9842 13398 9847 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 10374 13314 10402 13902
rect 10817 13846 10822 13874
rect 10850 13846 11326 13874
rect 11354 13846 11359 13874
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 10873 13454 10878 13482
rect 10906 13454 10911 13482
rect 10878 13426 10906 13454
rect 10878 13398 11998 13426
rect 12026 13398 12031 13426
rect 10369 13286 10374 13314
rect 10402 13286 10407 13314
rect 10878 13258 10906 13398
rect 7121 13230 7126 13258
rect 7154 13230 7630 13258
rect 7658 13230 7663 13258
rect 9529 13230 9534 13258
rect 9562 13230 9926 13258
rect 9954 13230 10906 13258
rect 6169 13174 6174 13202
rect 6202 13174 7742 13202
rect 7770 13174 7775 13202
rect 0 13146 400 13160
rect 0 13118 966 13146
rect 994 13118 999 13146
rect 2137 13118 2142 13146
rect 2170 13118 6062 13146
rect 6090 13118 7574 13146
rect 7602 13118 7607 13146
rect 8185 13118 8190 13146
rect 8218 13118 8694 13146
rect 8722 13118 8727 13146
rect 11545 13118 11550 13146
rect 11578 13118 11774 13146
rect 11802 13118 11807 13146
rect 11881 13118 11886 13146
rect 11914 13118 12614 13146
rect 12642 13118 12647 13146
rect 0 13104 400 13118
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 7345 12894 7350 12922
rect 7378 12894 7574 12922
rect 0 12810 400 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 0 12768 400 12782
rect 7546 12754 7574 12894
rect 7546 12726 7686 12754
rect 7714 12726 9086 12754
rect 9114 12726 9119 12754
rect 9249 12726 9254 12754
rect 9282 12726 9814 12754
rect 9842 12726 9847 12754
rect 7121 12670 7126 12698
rect 7154 12670 7462 12698
rect 7490 12670 7495 12698
rect 7546 12642 7574 12726
rect 7462 12614 7574 12642
rect 11545 12614 11550 12642
rect 11578 12614 13286 12642
rect 13314 12614 13319 12642
rect 7462 12586 7490 12614
rect 7457 12558 7462 12586
rect 7490 12558 7495 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 15946 12334 18830 12362
rect 18858 12334 18863 12362
rect 15946 12306 15974 12334
rect 7625 12278 7630 12306
rect 7658 12278 7854 12306
rect 7882 12278 8694 12306
rect 8722 12278 8918 12306
rect 8946 12278 10374 12306
rect 10402 12278 10710 12306
rect 10738 12278 11494 12306
rect 11522 12278 12166 12306
rect 12194 12278 12670 12306
rect 12698 12278 13006 12306
rect 13034 12278 13039 12306
rect 14065 12278 14070 12306
rect 14098 12278 14462 12306
rect 14490 12278 15974 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 13729 11998 13734 12026
rect 13762 11998 15974 12026
rect 15946 11970 15974 11998
rect 2137 11942 2142 11970
rect 2170 11942 4214 11970
rect 6897 11942 6902 11970
rect 6930 11942 7630 11970
rect 7658 11942 7663 11970
rect 15946 11942 18830 11970
rect 18858 11942 18863 11970
rect 4186 11914 4214 11942
rect 4186 11886 6958 11914
rect 6986 11886 6991 11914
rect 7905 11886 7910 11914
rect 7938 11886 8358 11914
rect 8386 11886 9926 11914
rect 9954 11886 10990 11914
rect 11018 11886 11023 11914
rect 12889 11886 12894 11914
rect 12922 11886 13902 11914
rect 13930 11886 13935 11914
rect 8017 11830 8022 11858
rect 8050 11830 8470 11858
rect 8498 11830 8503 11858
rect 9814 11830 9870 11858
rect 9898 11830 10122 11858
rect 11993 11830 11998 11858
rect 12026 11830 12278 11858
rect 12306 11830 12311 11858
rect 0 11802 400 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 0 11760 400 11774
rect 9814 11746 9842 11830
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 10094 11746 10122 11830
rect 20600 11802 21000 11816
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 20600 11760 21000 11774
rect 8689 11718 8694 11746
rect 8722 11718 9842 11746
rect 10094 11718 10458 11746
rect 11601 11718 11606 11746
rect 11634 11718 12054 11746
rect 12082 11718 12087 11746
rect 10430 11690 10458 11718
rect 9585 11662 9590 11690
rect 9618 11662 10318 11690
rect 10346 11662 10351 11690
rect 10430 11662 12502 11690
rect 12530 11662 12535 11690
rect 12777 11662 12782 11690
rect 12810 11662 13734 11690
rect 13762 11662 13767 11690
rect 8577 11606 8582 11634
rect 8610 11606 9030 11634
rect 9058 11606 9063 11634
rect 9641 11606 9646 11634
rect 9674 11606 11830 11634
rect 11858 11606 11863 11634
rect 12049 11606 12054 11634
rect 12082 11606 12838 11634
rect 12866 11606 12871 11634
rect 11046 11578 11074 11606
rect 2137 11550 2142 11578
rect 2170 11550 4214 11578
rect 8969 11550 8974 11578
rect 9002 11550 9310 11578
rect 9338 11550 9343 11578
rect 10201 11550 10206 11578
rect 10234 11550 10598 11578
rect 10626 11550 10631 11578
rect 11041 11550 11046 11578
rect 11074 11550 11079 11578
rect 4186 11522 4214 11550
rect 4186 11494 5334 11522
rect 5362 11494 5367 11522
rect 6953 11494 6958 11522
rect 6986 11494 8582 11522
rect 8610 11494 8615 11522
rect 10033 11494 10038 11522
rect 10066 11494 10262 11522
rect 10290 11494 11158 11522
rect 11186 11494 11191 11522
rect 0 11466 400 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 7401 11438 7406 11466
rect 7434 11438 7686 11466
rect 7714 11438 8862 11466
rect 8890 11438 8895 11466
rect 10873 11438 10878 11466
rect 10906 11438 11494 11466
rect 11522 11438 11527 11466
rect 0 11424 400 11438
rect 6953 11382 6958 11410
rect 6986 11382 8694 11410
rect 8722 11382 8727 11410
rect 10313 11382 10318 11410
rect 10346 11382 11102 11410
rect 11130 11382 11135 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9193 11326 9198 11354
rect 9226 11326 10710 11354
rect 10738 11326 12614 11354
rect 12642 11326 12647 11354
rect 7569 11270 7574 11298
rect 7602 11270 7966 11298
rect 7994 11270 9758 11298
rect 9786 11270 9791 11298
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 10145 11214 10150 11242
rect 10178 11214 10654 11242
rect 10682 11214 10687 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 2137 11158 2142 11186
rect 2170 11158 6622 11186
rect 6650 11158 6655 11186
rect 8801 11158 8806 11186
rect 8834 11158 8946 11186
rect 9025 11158 9030 11186
rect 9058 11158 10262 11186
rect 10290 11158 10295 11186
rect 8918 11130 8946 11158
rect 0 11102 994 11130
rect 6393 11102 6398 11130
rect 6426 11102 6734 11130
rect 6762 11102 6767 11130
rect 6897 11102 6902 11130
rect 6930 11102 7630 11130
rect 7658 11102 7663 11130
rect 8918 11102 8974 11130
rect 9002 11102 9007 11130
rect 0 11088 400 11102
rect 8801 11046 8806 11074
rect 8834 11046 9086 11074
rect 9114 11046 9119 11074
rect 5329 10990 5334 11018
rect 5362 10990 7630 11018
rect 7658 10990 7663 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 12273 10934 12278 10962
rect 12306 10934 12838 10962
rect 12866 10934 12871 10962
rect 6785 10878 6790 10906
rect 6818 10878 7126 10906
rect 7154 10878 7159 10906
rect 10537 10878 10542 10906
rect 10570 10878 12110 10906
rect 12138 10878 12894 10906
rect 12922 10878 13622 10906
rect 13650 10878 13655 10906
rect 9193 10822 9198 10850
rect 9226 10822 10374 10850
rect 10402 10822 10407 10850
rect 11937 10822 11942 10850
rect 11970 10822 12726 10850
rect 12754 10822 12759 10850
rect 0 10794 400 10808
rect 0 10766 994 10794
rect 2137 10766 2142 10794
rect 2170 10766 5222 10794
rect 5250 10766 5255 10794
rect 7961 10766 7966 10794
rect 7994 10766 8750 10794
rect 8778 10766 9142 10794
rect 9170 10766 9175 10794
rect 9697 10766 9702 10794
rect 9730 10766 9870 10794
rect 9898 10766 9903 10794
rect 0 10752 400 10766
rect 966 10738 994 10766
rect 961 10710 966 10738
rect 994 10710 999 10738
rect 6281 10710 6286 10738
rect 6314 10710 6902 10738
rect 6930 10710 6935 10738
rect 11209 10710 11214 10738
rect 11242 10710 11494 10738
rect 11522 10710 11527 10738
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 10929 10542 10934 10570
rect 10962 10542 11606 10570
rect 11634 10542 11639 10570
rect 8017 10430 8022 10458
rect 8050 10430 8638 10458
rect 8666 10430 9646 10458
rect 9674 10430 11214 10458
rect 11242 10430 11247 10458
rect 12553 10430 12558 10458
rect 12586 10430 14294 10458
rect 14322 10430 14327 10458
rect 5217 10374 5222 10402
rect 5250 10374 6902 10402
rect 6930 10374 7350 10402
rect 7378 10374 7383 10402
rect 9081 10374 9086 10402
rect 9114 10374 9870 10402
rect 9898 10374 9903 10402
rect 10313 10374 10318 10402
rect 10346 10374 10990 10402
rect 11018 10374 11774 10402
rect 11802 10374 12278 10402
rect 12306 10374 12311 10402
rect 2081 10262 2086 10290
rect 2114 10262 9478 10290
rect 9506 10262 9646 10290
rect 9674 10262 9679 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 7849 10094 7854 10122
rect 7882 10094 8526 10122
rect 8554 10094 8559 10122
rect 6337 10038 6342 10066
rect 6370 10038 6846 10066
rect 6874 10038 6879 10066
rect 8465 10038 8470 10066
rect 8498 10038 9198 10066
rect 9226 10038 9422 10066
rect 9450 10038 9455 10066
rect 9809 10038 9814 10066
rect 9842 10038 10934 10066
rect 10962 10038 10967 10066
rect 7401 9982 7406 10010
rect 7434 9982 8694 10010
rect 8722 9982 9030 10010
rect 9058 9982 9063 10010
rect 9137 9982 9142 10010
rect 9170 9982 11494 10010
rect 11522 9982 11527 10010
rect 15946 9982 18830 10010
rect 18858 9982 18863 10010
rect 9142 9954 9170 9982
rect 15946 9954 15974 9982
rect 8409 9926 8414 9954
rect 8442 9926 9170 9954
rect 12217 9926 12222 9954
rect 12250 9926 12614 9954
rect 12642 9926 12647 9954
rect 13953 9926 13958 9954
rect 13986 9926 14574 9954
rect 14602 9926 15974 9954
rect 6897 9870 6902 9898
rect 6930 9870 7966 9898
rect 7994 9870 7999 9898
rect 8129 9870 8134 9898
rect 8162 9870 8358 9898
rect 8386 9870 8391 9898
rect 9473 9870 9478 9898
rect 9506 9870 11886 9898
rect 11914 9870 13230 9898
rect 13258 9870 13263 9898
rect 8745 9814 8750 9842
rect 8778 9814 8862 9842
rect 8890 9814 10262 9842
rect 10290 9814 10295 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 10593 9758 10598 9786
rect 10626 9758 11102 9786
rect 11130 9758 11135 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 10201 9702 10206 9730
rect 10234 9702 10878 9730
rect 10906 9702 10911 9730
rect 11993 9702 11998 9730
rect 12026 9702 12502 9730
rect 12530 9702 12535 9730
rect 11321 9590 11326 9618
rect 11354 9590 11886 9618
rect 11914 9590 12222 9618
rect 12250 9590 12255 9618
rect 9249 9534 9254 9562
rect 9282 9534 10150 9562
rect 10178 9534 10183 9562
rect 12777 9534 12782 9562
rect 12810 9534 13342 9562
rect 13370 9534 13790 9562
rect 13818 9534 13823 9562
rect 7289 9478 7294 9506
rect 7322 9478 7742 9506
rect 7770 9478 8246 9506
rect 8274 9478 8279 9506
rect 8913 9478 8918 9506
rect 8946 9478 9310 9506
rect 9338 9478 9646 9506
rect 9674 9478 9679 9506
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 8577 9310 8582 9338
rect 8610 9310 8974 9338
rect 9002 9310 9814 9338
rect 9842 9310 10682 9338
rect 10817 9310 10822 9338
rect 10850 9310 11326 9338
rect 11354 9310 12054 9338
rect 12082 9310 12087 9338
rect 10654 9282 10682 9310
rect 9641 9254 9646 9282
rect 9674 9254 10094 9282
rect 10122 9254 10127 9282
rect 10649 9254 10654 9282
rect 10682 9254 10687 9282
rect 11153 9254 11158 9282
rect 11186 9254 11606 9282
rect 11634 9254 11639 9282
rect 6001 9198 6006 9226
rect 6034 9198 7518 9226
rect 7546 9198 7551 9226
rect 9025 9198 9030 9226
rect 9058 9198 9142 9226
rect 9170 9198 9366 9226
rect 9394 9198 9399 9226
rect 9529 9198 9534 9226
rect 9562 9198 9870 9226
rect 9898 9198 9903 9226
rect 11097 9198 11102 9226
rect 11130 9198 11438 9226
rect 11466 9198 12614 9226
rect 12642 9198 12647 9226
rect 9870 9170 9898 9198
rect 6393 9142 6398 9170
rect 6426 9142 7126 9170
rect 7154 9142 7159 9170
rect 9870 9142 11270 9170
rect 11298 9142 11303 9170
rect 7345 9030 7350 9058
rect 7378 9030 11438 9058
rect 11466 9030 11471 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 2137 8806 2142 8834
rect 2170 8806 5614 8834
rect 5642 8806 7182 8834
rect 7210 8806 7215 8834
rect 9585 8806 9590 8834
rect 9618 8806 9814 8834
rect 9842 8806 9847 8834
rect 11769 8806 11774 8834
rect 11802 8806 12054 8834
rect 12082 8806 12726 8834
rect 12754 8806 12759 8834
rect 0 8750 994 8778
rect 9310 8750 10262 8778
rect 10290 8750 10710 8778
rect 10738 8750 10743 8778
rect 0 8736 400 8750
rect 9310 8722 9338 8750
rect 7905 8694 7910 8722
rect 7938 8694 8358 8722
rect 8386 8694 9310 8722
rect 9338 8694 9343 8722
rect 9529 8694 9534 8722
rect 9562 8694 9870 8722
rect 9898 8694 10150 8722
rect 10178 8694 12278 8722
rect 12306 8694 13286 8722
rect 13314 8694 13319 8722
rect 8857 8638 8862 8666
rect 8890 8638 8946 8666
rect 8918 8442 8946 8638
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 20600 8442 21000 8456
rect 8913 8414 8918 8442
rect 8946 8414 8951 8442
rect 11377 8414 11382 8442
rect 11410 8414 12782 8442
rect 12810 8414 12815 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 20600 8400 21000 8414
rect 7009 8358 7014 8386
rect 7042 8358 7574 8386
rect 7602 8358 7607 8386
rect 10929 8358 10934 8386
rect 10962 8358 11662 8386
rect 11690 8358 11695 8386
rect 14401 8358 14406 8386
rect 14434 8358 18942 8386
rect 18970 8358 18975 8386
rect 8745 8302 8750 8330
rect 8778 8302 9030 8330
rect 9058 8302 11774 8330
rect 11802 8302 11807 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 13561 8190 13566 8218
rect 13594 8190 14406 8218
rect 14434 8190 14439 8218
rect 11153 8134 11158 8162
rect 11186 8134 12054 8162
rect 12082 8134 13174 8162
rect 13202 8134 13207 8162
rect 0 8106 400 8120
rect 20600 8106 21000 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 11601 8078 11606 8106
rect 11634 8078 12110 8106
rect 12138 8078 12950 8106
rect 12978 8078 12983 8106
rect 19945 8078 19950 8106
rect 19978 8078 21000 8106
rect 0 8064 400 8078
rect 20600 8064 21000 8078
rect 10089 8022 10094 8050
rect 10122 8022 10654 8050
rect 10682 8022 10687 8050
rect 11433 8022 11438 8050
rect 11466 8022 12502 8050
rect 12530 8022 12535 8050
rect 13057 8022 13062 8050
rect 13090 8022 13902 8050
rect 13930 8022 13935 8050
rect 10369 7966 10374 7994
rect 10402 7966 11158 7994
rect 11186 7966 11494 7994
rect 11522 7966 11830 7994
rect 11858 7966 11863 7994
rect 11937 7966 11942 7994
rect 11970 7966 12726 7994
rect 12754 7966 12759 7994
rect 7009 7910 7014 7938
rect 7042 7910 7574 7938
rect 10425 7910 10430 7938
rect 10458 7910 10878 7938
rect 10906 7910 10911 7938
rect 7546 7658 7574 7910
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 20600 7770 21000 7784
rect 9921 7742 9926 7770
rect 9954 7742 10766 7770
rect 10794 7742 10799 7770
rect 15946 7742 18830 7770
rect 18858 7742 18863 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 15946 7714 15974 7742
rect 20600 7728 21000 7742
rect 14849 7686 14854 7714
rect 14882 7686 15974 7714
rect 7546 7630 8750 7658
rect 8778 7630 9758 7658
rect 9786 7630 10038 7658
rect 10066 7630 10071 7658
rect 14009 7630 14014 7658
rect 14042 7630 14742 7658
rect 14770 7630 18774 7658
rect 18802 7630 18807 7658
rect 2137 7574 2142 7602
rect 2170 7574 5894 7602
rect 5922 7574 6846 7602
rect 6874 7574 6879 7602
rect 7569 7574 7574 7602
rect 7602 7574 9198 7602
rect 9226 7574 9231 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 20600 7434 21000 7448
rect 20001 7406 20006 7434
rect 20034 7406 21000 7434
rect 20600 7392 21000 7406
rect 8913 7294 8918 7322
rect 8946 7294 9198 7322
rect 9226 7294 10794 7322
rect 10766 7266 10794 7294
rect 10761 7238 10766 7266
rect 10794 7238 11326 7266
rect 11354 7238 11774 7266
rect 11802 7238 11807 7266
rect 14737 7126 14742 7154
rect 14770 7126 18830 7154
rect 18858 7126 18863 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 10145 6846 10150 6874
rect 10178 6846 10766 6874
rect 10794 6846 10799 6874
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9809 6510 9814 6538
rect 9842 6510 10318 6538
rect 10346 6510 10351 6538
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 12777 2030 12782 2058
rect 12810 2030 13398 2058
rect 13426 2030 13431 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 12441 1806 12446 1834
rect 12474 1806 13062 1834
rect 13090 1806 13095 1834
rect 10089 1694 10094 1722
rect 10122 1694 10878 1722
rect 10906 1694 10911 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12768 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11536 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11536 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10024 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12656 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _106_
timestamp 1698175906
transform -1 0 11200 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _107_
timestamp 1698175906
transform 1 0 10136 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _108_
timestamp 1698175906
transform -1 0 8960 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform 1 0 9576 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9128 0 -1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _113_
timestamp 1698175906
transform -1 0 8512 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _114_
timestamp 1698175906
transform 1 0 12432 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform -1 0 11872 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_
timestamp 1698175906
transform -1 0 11424 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 11424 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _118_
timestamp 1698175906
transform -1 0 12600 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 12544 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9128 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _121_
timestamp 1698175906
transform -1 0 8960 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_
timestamp 1698175906
transform -1 0 9968 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10136 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 8624 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11312 0 1 8624
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _128_
timestamp 1698175906
transform -1 0 13776 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698175906
transform -1 0 13496 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _130_
timestamp 1698175906
transform 1 0 9128 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_
timestamp 1698175906
transform -1 0 8680 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _132_
timestamp 1698175906
transform -1 0 8232 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_
timestamp 1698175906
transform -1 0 7000 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12152 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11368 0 -1 10976
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _136_
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _137_
timestamp 1698175906
transform 1 0 12992 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform 1 0 10024 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform 1 0 10192 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _140_
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _141_
timestamp 1698175906
transform 1 0 8960 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11368 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform -1 0 9520 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform 1 0 9688 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 10976 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 10472 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9128 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _148_
timestamp 1698175906
transform 1 0 13720 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform -1 0 12376 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13160 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _151_
timestamp 1698175906
transform -1 0 11648 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform 1 0 8680 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform -1 0 9632 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 9128 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _155_
timestamp 1698175906
transform 1 0 13776 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _156_
timestamp 1698175906
transform -1 0 12208 0 1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12880 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform 1 0 8792 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 1051 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform -1 0 8512 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _161_
timestamp 1698175906
transform 1 0 7560 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform 1 0 9800 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _163_
timestamp 1698175906
transform 1 0 9800 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _164_
timestamp 1698175906
transform -1 0 9352 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _165_
timestamp 1698175906
transform 1 0 10136 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10024 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _167_
timestamp 1698175906
transform -1 0 10136 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8120 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _169_
timestamp 1698175906
transform -1 0 7000 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 7112 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform 1 0 7168 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _172_
timestamp 1698175906
transform 1 0 11760 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform 1 0 11592 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _174_
timestamp 1698175906
transform -1 0 9632 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _175_
timestamp 1698175906
transform 1 0 9128 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform 1 0 9744 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _177_
timestamp 1698175906
transform 1 0 9240 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11424 0 1 10192
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _179_
timestamp 1698175906
transform 1 0 7000 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _181_
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _182_
timestamp 1698175906
transform -1 0 9352 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _183_
timestamp 1698175906
transform 1 0 8512 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _184_
timestamp 1698175906
transform 1 0 8344 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _186_
timestamp 1698175906
transform 1 0 13832 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _187_
timestamp 1698175906
transform -1 0 13552 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform -1 0 7504 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _189_
timestamp 1698175906
transform 1 0 6776 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform -1 0 7728 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7224 0 1 12544
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _192_
timestamp 1698175906
transform -1 0 10472 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1698175906
transform 1 0 11368 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _194_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 -1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _195_
timestamp 1698175906
transform -1 0 12768 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 1331 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _197_
timestamp 1698175906
transform 1 0 11592 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _198_
timestamp 1698175906
transform -1 0 12992 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _199_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 -1 11760
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_
timestamp 1698175906
transform -1 0 7896 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _201_
timestamp 1698175906
transform -1 0 7448 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7504 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 8792 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 12880 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 7448 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 5880 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 12768 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 10024 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 9800 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 13048 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 8120 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 12992 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 6888 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform -1 0 7448 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 11200 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform -1 0 7168 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 8512 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 12936 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform -1 0 6776 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform -1 0 7616 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 11368 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 12208 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 7728 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _228_
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _229_
timestamp 1698175906
transform -1 0 7000 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _230_
timestamp 1698175906
transform 1 0 12824 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _231_
timestamp 1698175906
transform 1 0 14616 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform -1 0 10808 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 12768 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 9184 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform -1 0 7728 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform -1 0 12992 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 11760 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 11536 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 12936 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform -1 0 9856 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 12880 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 6888 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 7560 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 13272 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 10360 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 7560 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 8904 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 7112 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 8008 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 12096 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 7840 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9576 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 9576 0 -1 8624
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 9520 0 -1 12544
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 11760 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 11984 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12432 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 13944 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 12208 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 12768 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 14280 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 16072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 16296 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 8456 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1698175906
transform 1 0 8680 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_181
timestamp 1698175906
transform 1 0 10808 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_166
timestamp 1698175906
transform 1 0 9968 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_196
timestamp 1698175906
transform 1 0 11648 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_200
timestamp 1698175906
transform 1 0 11872 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698175906
transform 1 0 7336 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_121
timestamp 1698175906
transform 1 0 7448 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_151
timestamp 1698175906
transform 1 0 9128 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_155
timestamp 1698175906
transform 1 0 9352 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_159
timestamp 1698175906
transform 1 0 9576 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_166
timestamp 1698175906
transform 1 0 9968 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 10416 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_185
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_187
timestamp 1698175906
transform 1 0 11144 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_223
timestamp 1698175906
transform 1 0 13160 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_227
timestamp 1698175906
transform 1 0 13384 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 14280 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_253
timestamp 1698175906
transform 1 0 14840 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_285
timestamp 1698175906
transform 1 0 16632 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_301
timestamp 1698175906
transform 1 0 17528 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_309
timestamp 1698175906
transform 1 0 17976 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_313
timestamp 1698175906
transform 1 0 18200 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698175906
transform 1 0 5600 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_121
timestamp 1698175906
transform 1 0 7448 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_125
timestamp 1698175906
transform 1 0 7672 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698175906
transform 1 0 8120 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698175906
transform 1 0 8344 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 8456 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_151
timestamp 1698175906
transform 1 0 9128 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_159
timestamp 1698175906
transform 1 0 9576 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_169
timestamp 1698175906
transform 1 0 10136 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_185
timestamp 1698175906
transform 1 0 11032 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_193
timestamp 1698175906
transform 1 0 11480 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698175906
transform 1 0 12040 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 12264 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698175906
transform 1 0 12768 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_255
timestamp 1698175906
transform 1 0 14952 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_271
timestamp 1698175906
transform 1 0 15848 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 18704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_109
timestamp 1698175906
transform 1 0 6776 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698175906
transform 1 0 7336 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_150
timestamp 1698175906
transform 1 0 9072 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_154
timestamp 1698175906
transform 1 0 9296 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_185
timestamp 1698175906
transform 1 0 11032 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_208
timestamp 1698175906
transform 1 0 12320 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698175906
transform 1 0 14112 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 5152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_84
timestamp 1698175906
transform 1 0 5376 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_86
timestamp 1698175906
transform 1 0 5488 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_121
timestamp 1698175906
transform 1 0 7448 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_125
timestamp 1698175906
transform 1 0 7672 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698175906
transform 1 0 8120 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 8344 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_148
timestamp 1698175906
transform 1 0 8960 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_156
timestamp 1698175906
transform 1 0 9408 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_158
timestamp 1698175906
transform 1 0 9520 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_247
timestamp 1698175906
transform 1 0 14504 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_131
timestamp 1698175906
transform 1 0 8008 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_135
timestamp 1698175906
transform 1 0 8232 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_152
timestamp 1698175906
transform 1 0 9184 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_160
timestamp 1698175906
transform 1 0 9632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_212
timestamp 1698175906
transform 1 0 12544 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_220
timestamp 1698175906
transform 1 0 12992 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_222
timestamp 1698175906
transform 1 0 13104 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_229
timestamp 1698175906
transform 1 0 13496 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_104
timestamp 1698175906
transform 1 0 6496 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_112
timestamp 1698175906
transform 1 0 6944 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_121
timestamp 1698175906
transform 1 0 7448 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698175906
transform 1 0 8344 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_159
timestamp 1698175906
transform 1 0 9576 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_172
timestamp 1698175906
transform 1 0 10304 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_200
timestamp 1698175906
transform 1 0 11872 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_218
timestamp 1698175906
transform 1 0 12880 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_250
timestamp 1698175906
transform 1 0 14672 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_266
timestamp 1698175906
transform 1 0 15568 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 16016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_113
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_129
timestamp 1698175906
transform 1 0 7896 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_165
timestamp 1698175906
transform 1 0 9912 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698175906
transform 1 0 11032 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_213
timestamp 1698175906
transform 1 0 12600 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_217
timestamp 1698175906
transform 1 0 12824 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_221
timestamp 1698175906
transform 1 0 13048 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_239
timestamp 1698175906
transform 1 0 14056 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 14280 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_92
timestamp 1698175906
transform 1 0 5824 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_122
timestamp 1698175906
transform 1 0 7504 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_126
timestamp 1698175906
transform 1 0 7728 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_128
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_148
timestamp 1698175906
transform 1 0 8960 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698175906
transform 1 0 9072 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_216
timestamp 1698175906
transform 1 0 12768 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_220
timestamp 1698175906
transform 1 0 12992 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_250
timestamp 1698175906
transform 1 0 14672 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_266
timestamp 1698175906
transform 1 0 15568 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_113
timestamp 1698175906
transform 1 0 7000 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_117
timestamp 1698175906
transform 1 0 7224 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_133
timestamp 1698175906
transform 1 0 8120 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_137
timestamp 1698175906
transform 1 0 8344 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_139
timestamp 1698175906
transform 1 0 8456 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_152
timestamp 1698175906
transform 1 0 9184 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_156
timestamp 1698175906
transform 1 0 9408 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_159
timestamp 1698175906
transform 1 0 9576 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_169
timestamp 1698175906
transform 1 0 10136 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 10360 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_214
timestamp 1698175906
transform 1 0 12656 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_122
timestamp 1698175906
transform 1 0 7504 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_132
timestamp 1698175906
transform 1 0 8064 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_148
timestamp 1698175906
transform 1 0 8960 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_155
timestamp 1698175906
transform 1 0 9352 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_226
timestamp 1698175906
transform 1 0 13328 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_258
timestamp 1698175906
transform 1 0 15120 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 16016 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_113
timestamp 1698175906
transform 1 0 7000 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_121
timestamp 1698175906
transform 1 0 7448 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_133
timestamp 1698175906
transform 1 0 8120 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_137
timestamp 1698175906
transform 1 0 8344 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_139
timestamp 1698175906
transform 1 0 8456 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_155
timestamp 1698175906
transform 1 0 9352 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_163
timestamp 1698175906
transform 1 0 9800 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_200
timestamp 1698175906
transform 1 0 11872 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_206
timestamp 1698175906
transform 1 0 12208 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_238
timestamp 1698175906
transform 1 0 14000 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 14224 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_80
timestamp 1698175906
transform 1 0 5152 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_160
timestamp 1698175906
transform 1 0 9632 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_188
timestamp 1698175906
transform 1 0 11200 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_190
timestamp 1698175906
transform 1 0 11312 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_197
timestamp 1698175906
transform 1 0 11704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_220
timestamp 1698175906
transform 1 0 12992 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_252
timestamp 1698175906
transform 1 0 14784 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_268
timestamp 1698175906
transform 1 0 15680 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_113
timestamp 1698175906
transform 1 0 7000 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_129
timestamp 1698175906
transform 1 0 7896 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_145
timestamp 1698175906
transform 1 0 8792 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_149
timestamp 1698175906
transform 1 0 9016 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_157
timestamp 1698175906
transform 1 0 9464 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_161
timestamp 1698175906
transform 1 0 9688 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_169
timestamp 1698175906
transform 1 0 10136 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 10360 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_96
timestamp 1698175906
transform 1 0 6048 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_126
timestamp 1698175906
transform 1 0 7728 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698175906
transform 1 0 7952 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 12320 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_216
timestamp 1698175906
transform 1 0 12768 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_218
timestamp 1698175906
transform 1 0 12880 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_248
timestamp 1698175906
transform 1 0 14560 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_128
timestamp 1698175906
transform 1 0 7840 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_144
timestamp 1698175906
transform 1 0 8736 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_152
timestamp 1698175906
transform 1 0 9184 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_167
timestamp 1698175906
transform 1 0 10024 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_220
timestamp 1698175906
transform 1 0 12992 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_230
timestamp 1698175906
transform 1 0 13552 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 14000 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_92
timestamp 1698175906
transform 1 0 5824 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_94
timestamp 1698175906
transform 1 0 5936 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_129
timestamp 1698175906
transform 1 0 7896 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698175906
transform 1 0 8120 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698175906
transform 1 0 8344 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_171
timestamp 1698175906
transform 1 0 10248 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_175
timestamp 1698175906
transform 1 0 10472 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_191
timestamp 1698175906
transform 1 0 11368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_204
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_216
timestamp 1698175906
transform 1 0 12768 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 2240 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 2464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_126
timestamp 1698175906
transform 1 0 7728 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_130
timestamp 1698175906
transform 1 0 7952 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_132
timestamp 1698175906
transform 1 0 8064 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_167
timestamp 1698175906
transform 1 0 10024 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_169
timestamp 1698175906
transform 1 0 10136 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_184
timestamp 1698175906
transform 1 0 10976 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_216
timestamp 1698175906
transform 1 0 12768 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_232
timestamp 1698175906
transform 1 0 13664 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_240
timestamp 1698175906
transform 1 0 14112 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_151
timestamp 1698175906
transform 1 0 9128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_160
timestamp 1698175906
transform 1 0 9632 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_162
timestamp 1698175906
transform 1 0 9744 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_192
timestamp 1698175906
transform 1 0 11424 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_196
timestamp 1698175906
transform 1 0 11648 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 12320 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_139
timestamp 1698175906
transform 1 0 8456 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_155
timestamp 1698175906
transform 1 0 9352 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_159
timestamp 1698175906
transform 1 0 9576 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_161
timestamp 1698175906
transform 1 0 9688 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_164
timestamp 1698175906
transform 1 0 9856 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 10304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 10416 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_158
timestamp 1698175906
transform 1 0 9520 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_166
timestamp 1698175906
transform 1 0 9968 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 10080 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 11592 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 12040 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 14280 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 16072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_245
timestamp 1698175906
transform 1 0 14392 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_261
timestamp 1698175906
transform 1 0 15288 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_269
timestamp 1698175906
transform 1 0 15736 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698175906
transform 1 0 15848 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita61_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12432 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita61_26
timestamp 1698175906
transform -1 0 14392 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 12824 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 10136 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 12824 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 12488 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 12096 0 12152 400 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 7392 21000 7448 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 14112 20600 14168 21000 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 10752 400 10808 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 12768 0 12824 400 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 13468 9716 13468 9716 0 _000_
rlabel metal2 8596 13748 8596 13748 0 _001_
rlabel metal2 13300 7840 13300 7840 0 _002_
rlabel metal3 6580 11116 6580 11116 0 _003_
rlabel metal2 6972 7756 6972 7756 0 _004_
rlabel metal2 11676 7434 11676 7434 0 _005_
rlabel metal2 9380 12936 9380 12936 0 _006_
rlabel metal2 6468 8260 6468 8260 0 _007_
rlabel metal2 8036 11732 8036 11732 0 _008_
rlabel metal2 13412 12516 13412 12516 0 _009_
rlabel metal3 6608 10724 6608 10724 0 _010_
rlabel metal3 7308 12684 7308 12684 0 _011_
rlabel metal2 11060 11788 11060 11788 0 _012_
rlabel metal2 11844 12936 11844 12936 0 _013_
rlabel metal2 12348 11704 12348 11704 0 _014_
rlabel metal2 7252 12600 7252 12600 0 _015_
rlabel metal2 8372 7084 8372 7084 0 _016_
rlabel metal2 9296 6524 9296 6524 0 _017_
rlabel metal2 13356 8596 13356 8596 0 _018_
rlabel metal3 8148 8708 8148 8708 0 _019_
rlabel metal3 6608 10052 6608 10052 0 _020_
rlabel metal2 13244 10640 13244 10640 0 _021_
rlabel metal2 10500 7168 10500 7168 0 _022_
rlabel metal2 10304 13636 10304 13636 0 _023_
rlabel metal3 9156 11564 9156 11564 0 _024_
rlabel metal3 9212 13916 9212 13916 0 _025_
rlabel metal3 13496 8036 13496 8036 0 _026_
rlabel metal2 11620 8204 11620 8204 0 _027_
rlabel metal2 8820 11368 8820 11368 0 _028_
rlabel metal2 7420 12068 7420 12068 0 _029_
rlabel metal2 7308 9016 7308 9016 0 _030_
rlabel metal2 7812 11032 7812 11032 0 _031_
rlabel metal2 10108 11004 10108 11004 0 _032_
rlabel metal2 8400 11956 8400 11956 0 _033_
rlabel metal2 9072 10892 9072 10892 0 _034_
rlabel metal3 10724 11508 10724 11508 0 _035_
rlabel metal2 10080 11228 10080 11228 0 _036_
rlabel metal3 7784 11284 7784 11284 0 _037_
rlabel metal3 7280 11116 7280 11116 0 _038_
rlabel metal2 6972 8176 6972 8176 0 _039_
rlabel metal2 11900 7784 11900 7784 0 _040_
rlabel metal2 9492 9044 9492 9044 0 _041_
rlabel metal2 9352 9324 9352 9324 0 _042_
rlabel metal2 9800 13636 9800 13636 0 _043_
rlabel metal2 7364 9128 7364 9128 0 _044_
rlabel metal2 6412 8624 6412 8624 0 _045_
rlabel metal2 9212 11256 9212 11256 0 _046_
rlabel metal2 7364 13160 7364 13160 0 _047_
rlabel metal2 8764 11564 8764 11564 0 _048_
rlabel metal2 11452 11424 11452 11424 0 _049_
rlabel metal2 13972 12348 13972 12348 0 _050_
rlabel metal2 7252 10808 7252 10808 0 _051_
rlabel metal2 7336 12684 7336 12684 0 _052_
rlabel metal2 10332 9072 10332 9072 0 _053_
rlabel metal2 11508 11480 11508 11480 0 _054_
rlabel metal3 12264 13132 12264 13132 0 _055_
rlabel metal2 11676 12180 11676 12180 0 _056_
rlabel metal3 12460 11620 12460 11620 0 _057_
rlabel metal2 7140 13328 7140 13328 0 _058_
rlabel metal3 12432 9940 12432 9940 0 _059_
rlabel metal3 12040 9212 12040 9212 0 _060_
rlabel metal3 9716 9212 9716 9212 0 _061_
rlabel metal2 9968 7196 9968 7196 0 _062_
rlabel metal3 10668 10388 10668 10388 0 _063_
rlabel metal2 10948 10696 10948 10696 0 _064_
rlabel metal2 10276 9744 10276 9744 0 _065_
rlabel metal2 8680 8820 8680 8820 0 _066_
rlabel metal2 9660 9380 9660 9380 0 _067_
rlabel metal2 9828 9408 9828 9408 0 _068_
rlabel metal2 11788 8008 11788 8008 0 _069_
rlabel metal2 8652 7756 8652 7756 0 _070_
rlabel metal3 12404 8820 12404 8820 0 _071_
rlabel metal2 10556 10388 10556 10388 0 _072_
rlabel metal2 10360 7980 10360 7980 0 _073_
rlabel metal2 11844 11592 11844 11592 0 _074_
rlabel metal2 11312 9604 11312 9604 0 _075_
rlabel metal3 12796 8708 12796 8708 0 _076_
rlabel metal2 8820 10052 8820 10052 0 _077_
rlabel metal2 11228 10584 11228 10584 0 _078_
rlabel metal2 10080 7756 10080 7756 0 _079_
rlabel metal2 9828 7532 9828 7532 0 _080_
rlabel metal3 11620 8148 11620 8148 0 _081_
rlabel metal2 13776 8036 13776 8036 0 _082_
rlabel metal2 13636 8204 13636 8204 0 _083_
rlabel metal2 9212 10808 9212 10808 0 _084_
rlabel via2 8372 9884 8372 9884 0 _085_
rlabel metal2 6916 9744 6916 9744 0 _086_
rlabel metal2 6972 11144 6972 11144 0 _087_
rlabel metal2 11956 11144 11956 11144 0 _088_
rlabel metal2 12992 10780 12992 10780 0 _089_
rlabel metal2 10332 9324 10332 9324 0 _090_
rlabel metal3 10668 7924 10668 7924 0 _091_
rlabel metal2 9884 10584 9884 10584 0 _092_
rlabel metal2 9576 11564 9576 11564 0 _093_
rlabel metal2 7728 13468 7728 13468 0 _094_
rlabel metal2 12012 12488 12012 12488 0 _095_
rlabel metal2 10556 13468 10556 13468 0 _096_
rlabel metal2 11900 10164 11900 10164 0 _097_
rlabel metal2 13524 9604 13524 9604 0 _098_
rlabel metal2 13636 10248 13636 10248 0 _099_
rlabel metal2 11564 10780 11564 10780 0 _100_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal3 10388 10052 10388 10052 0 clknet_0_clk
rlabel metal2 11788 7112 11788 7112 0 clknet_1_0__leaf_clk
rlabel metal2 6804 11760 6804 11760 0 clknet_1_1__leaf_clk
rlabel metal2 9268 9576 9268 9576 0 dut61.count\[0\]
rlabel metal2 7420 9968 7420 9968 0 dut61.count\[1\]
rlabel metal2 12572 10416 12572 10416 0 dut61.count\[2\]
rlabel metal2 11564 7182 11564 7182 0 dut61.count\[3\]
rlabel metal2 12208 15960 12208 15960 0 net1
rlabel metal2 6076 13104 6076 13104 0 net10
rlabel metal2 12908 3178 12908 3178 0 net11
rlabel metal2 12628 2982 12628 2982 0 net12
rlabel metal2 2156 8008 2156 8008 0 net13
rlabel metal3 3178 11956 3178 11956 0 net14
rlabel metal2 14084 12124 14084 12124 0 net15
rlabel metal3 3178 11564 3178 11564 0 net16
rlabel metal3 15414 7700 15414 7700 0 net17
rlabel metal2 9660 13804 9660 13804 0 net18
rlabel metal2 13972 9772 13972 9772 0 net19
rlabel metal2 12796 15960 12796 15960 0 net2
rlabel metal3 11088 13860 11088 13860 0 net20
rlabel metal2 13580 8120 13580 8120 0 net21
rlabel metal2 10388 2982 10388 2982 0 net22
rlabel metal2 5628 8596 5628 8596 0 net23
rlabel metal2 8820 2982 8820 2982 0 net24
rlabel metal2 12124 1015 12124 1015 0 net25
rlabel metal2 14196 18956 14196 18956 0 net26
rlabel metal2 13748 11844 13748 11844 0 net3
rlabel metal2 6188 12908 6188 12908 0 net4
rlabel metal2 18844 7392 18844 7392 0 net5
rlabel metal2 6748 10500 6748 10500 0 net6
rlabel metal2 14532 7616 14532 7616 0 net7
rlabel metal2 5236 10752 5236 10752 0 net8
rlabel metal2 10192 13524 10192 13524 0 net9
rlabel metal2 11788 19873 11788 19873 0 segm[10]
rlabel metal2 12796 19957 12796 19957 0 segm[11]
rlabel metal2 20020 11900 20020 11900 0 segm[12]
rlabel metal3 679 13132 679 13132 0 segm[13]
rlabel metal2 20020 7504 20020 7504 0 segm[1]
rlabel metal3 679 11116 679 11116 0 segm[2]
rlabel metal2 19964 8232 19964 8232 0 segm[4]
rlabel metal3 679 10780 679 10780 0 segm[5]
rlabel metal2 10108 19677 10108 19677 0 segm[6]
rlabel metal3 679 12796 679 12796 0 segm[7]
rlabel metal2 12796 1211 12796 1211 0 segm[8]
rlabel metal2 12460 1099 12460 1099 0 segm[9]
rlabel metal3 679 8092 679 8092 0 sel[0]
rlabel metal3 679 11788 679 11788 0 sel[10]
rlabel metal2 20020 12180 20020 12180 0 sel[11]
rlabel metal3 679 11452 679 11452 0 sel[1]
rlabel metal2 20020 7924 20020 7924 0 sel[2]
rlabel metal2 9436 19845 9436 19845 0 sel[3]
rlabel metal2 20020 9828 20020 9828 0 sel[4]
rlabel metal2 11116 19873 11116 19873 0 sel[5]
rlabel metal2 20020 8652 20020 8652 0 sel[6]
rlabel metal2 10108 1043 10108 1043 0 sel[7]
rlabel metal3 679 8764 679 8764 0 sel[8]
rlabel metal2 9100 1099 9100 1099 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
