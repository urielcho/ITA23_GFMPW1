magic
tech gf180mcuD
magscale 1 5
timestamp 1699643937
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11047 19137 11073 19143
rect 11047 19105 11073 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 8801 18999 8807 19025
rect 8833 18999 8839 19025
rect 10537 18999 10543 19025
rect 10569 18999 10575 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9199 18745 9225 18751
rect 9199 18713 9225 18719
rect 10151 18745 10177 18751
rect 10151 18713 10177 18719
rect 13399 18745 13425 18751
rect 13399 18713 13425 18719
rect 8801 18607 8807 18633
rect 8833 18607 8839 18633
rect 12889 18607 12895 18633
rect 12921 18607 12927 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 20119 17345 20145 17351
rect 20119 17313 20145 17319
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 8521 14351 8527 14377
rect 8553 14351 8559 14377
rect 12105 14351 12111 14377
rect 12137 14351 12143 14377
rect 12335 14321 12361 14327
rect 7121 14295 7127 14321
rect 7153 14295 7159 14321
rect 10705 14295 10711 14321
rect 10737 14295 10743 14321
rect 11041 14295 11047 14321
rect 11073 14295 11079 14321
rect 12335 14289 12361 14295
rect 7457 14239 7463 14265
rect 7489 14239 7495 14265
rect 8863 14209 8889 14215
rect 8863 14177 8889 14183
rect 9087 14209 9113 14215
rect 9087 14177 9113 14183
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8191 14041 8217 14047
rect 8191 14009 8217 14015
rect 10879 14041 10905 14047
rect 10879 14009 10905 14015
rect 8751 13985 8777 13991
rect 8751 13953 8777 13959
rect 10711 13985 10737 13991
rect 10711 13953 10737 13959
rect 11271 13985 11297 13991
rect 11271 13953 11297 13959
rect 8135 13929 8161 13935
rect 8135 13897 8161 13903
rect 8247 13929 8273 13935
rect 8247 13897 8273 13903
rect 8471 13929 8497 13935
rect 8471 13897 8497 13903
rect 8695 13929 8721 13935
rect 10823 13929 10849 13935
rect 9025 13903 9031 13929
rect 9057 13903 9063 13929
rect 8695 13897 8721 13903
rect 10823 13897 10849 13903
rect 10935 13929 10961 13935
rect 10935 13897 10961 13903
rect 11215 13929 11241 13935
rect 11215 13897 11241 13903
rect 9417 13847 9423 13873
rect 9449 13847 9455 13873
rect 10481 13847 10487 13873
rect 10513 13847 10519 13873
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 9199 13593 9225 13599
rect 8521 13567 8527 13593
rect 8553 13567 8559 13593
rect 9529 13567 9535 13593
rect 9561 13567 9567 13593
rect 12889 13567 12895 13593
rect 12921 13567 12927 13593
rect 9199 13561 9225 13567
rect 8807 13537 8833 13543
rect 7121 13511 7127 13537
rect 7153 13511 7159 13537
rect 8807 13505 8833 13511
rect 8919 13537 8945 13543
rect 9591 13537 9617 13543
rect 10095 13537 10121 13543
rect 9473 13511 9479 13537
rect 9505 13511 9511 13537
rect 9809 13511 9815 13537
rect 9841 13511 9847 13537
rect 8919 13505 8945 13511
rect 9591 13505 9617 13511
rect 10095 13505 10121 13511
rect 10375 13537 10401 13543
rect 11433 13511 11439 13537
rect 11465 13511 11471 13537
rect 10375 13505 10401 13511
rect 8695 13481 8721 13487
rect 7457 13455 7463 13481
rect 7489 13455 7495 13481
rect 8695 13449 8721 13455
rect 8751 13481 8777 13487
rect 8751 13449 8777 13455
rect 10151 13481 10177 13487
rect 11825 13455 11831 13481
rect 11857 13455 11863 13481
rect 10151 13449 10177 13455
rect 9703 13425 9729 13431
rect 9703 13393 9729 13399
rect 10039 13425 10065 13431
rect 10039 13393 10065 13399
rect 13119 13425 13145 13431
rect 13119 13393 13145 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8863 13257 8889 13263
rect 11607 13257 11633 13263
rect 10873 13231 10879 13257
rect 10905 13231 10911 13257
rect 8863 13225 8889 13231
rect 11607 13225 11633 13231
rect 8695 13201 8721 13207
rect 8695 13169 8721 13175
rect 12671 13201 12697 13207
rect 12671 13169 12697 13175
rect 8807 13145 8833 13151
rect 8807 13113 8833 13119
rect 8919 13145 8945 13151
rect 8919 13113 8945 13119
rect 8975 13145 9001 13151
rect 8975 13113 9001 13119
rect 11047 13145 11073 13151
rect 11047 13113 11073 13119
rect 11551 13145 11577 13151
rect 11551 13113 11577 13119
rect 11663 13145 11689 13151
rect 11663 13113 11689 13119
rect 12615 13145 12641 13151
rect 12615 13113 12641 13119
rect 11439 13089 11465 13095
rect 11439 13057 11465 13063
rect 11215 13033 11241 13039
rect 11215 13001 11241 13007
rect 11327 13033 11353 13039
rect 11327 13001 11353 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 8135 12865 8161 12871
rect 8135 12833 8161 12839
rect 9927 12865 9953 12871
rect 9927 12833 9953 12839
rect 10711 12865 10737 12871
rect 10711 12833 10737 12839
rect 9031 12809 9057 12815
rect 12671 12809 12697 12815
rect 12441 12783 12447 12809
rect 12473 12783 12479 12809
rect 9031 12777 9057 12783
rect 12671 12777 12697 12783
rect 8191 12753 8217 12759
rect 10985 12727 10991 12753
rect 11017 12727 11023 12753
rect 8191 12721 8217 12727
rect 8919 12697 8945 12703
rect 8919 12665 8945 12671
rect 9871 12697 9897 12703
rect 9871 12665 9897 12671
rect 10655 12697 10681 12703
rect 11377 12671 11383 12697
rect 11409 12671 11415 12697
rect 10655 12665 10681 12671
rect 7911 12641 7937 12647
rect 7911 12609 7937 12615
rect 8135 12641 8161 12647
rect 8527 12641 8553 12647
rect 8353 12615 8359 12641
rect 8385 12615 8391 12641
rect 8135 12609 8161 12615
rect 8527 12609 8553 12615
rect 8975 12641 9001 12647
rect 8975 12609 9001 12615
rect 9927 12641 9953 12647
rect 9927 12609 9953 12615
rect 10711 12641 10737 12647
rect 10711 12609 10737 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 8863 12473 8889 12479
rect 8863 12441 8889 12447
rect 11663 12473 11689 12479
rect 11663 12441 11689 12447
rect 12111 12473 12137 12479
rect 12111 12441 12137 12447
rect 8247 12417 8273 12423
rect 8247 12385 8273 12391
rect 8919 12417 8945 12423
rect 10257 12391 10263 12417
rect 10289 12391 10295 12417
rect 8919 12385 8945 12391
rect 9647 12361 9673 12367
rect 6449 12335 6455 12361
rect 6481 12335 6487 12361
rect 8353 12335 8359 12361
rect 8385 12335 8391 12361
rect 10145 12335 10151 12361
rect 10177 12335 10183 12361
rect 9647 12329 9673 12335
rect 11383 12305 11409 12311
rect 6841 12279 6847 12305
rect 6873 12279 6879 12305
rect 7905 12279 7911 12305
rect 7937 12279 7943 12305
rect 9417 12279 9423 12305
rect 9449 12279 9455 12305
rect 11881 12279 11887 12305
rect 11913 12279 11919 12305
rect 11383 12273 11409 12279
rect 8807 12249 8833 12255
rect 8807 12217 8833 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 967 12025 993 12031
rect 8191 12025 8217 12031
rect 4993 11999 4999 12025
rect 5025 11999 5031 12025
rect 967 11993 993 11999
rect 8191 11993 8217 11999
rect 8415 12025 8441 12031
rect 8415 11993 8441 11999
rect 9591 12025 9617 12031
rect 9591 11993 9617 11999
rect 10655 12025 10681 12031
rect 20007 12025 20033 12031
rect 13057 11999 13063 12025
rect 13089 11999 13095 12025
rect 10655 11993 10681 11999
rect 20007 11993 20033 11999
rect 7855 11969 7881 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 6393 11943 6399 11969
rect 6425 11943 6431 11969
rect 7855 11937 7881 11943
rect 8303 11969 8329 11975
rect 8303 11937 8329 11943
rect 8527 11969 8553 11975
rect 9361 11943 9367 11969
rect 9393 11943 9399 11969
rect 9977 11943 9983 11969
rect 10009 11943 10015 11969
rect 11041 11943 11047 11969
rect 11073 11943 11079 11969
rect 13953 11943 13959 11969
rect 13985 11943 13991 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 8527 11937 8553 11943
rect 12895 11913 12921 11919
rect 6057 11887 6063 11913
rect 6089 11887 6095 11913
rect 8577 11887 8583 11913
rect 8609 11887 8615 11913
rect 8969 11887 8975 11913
rect 9001 11887 9007 11913
rect 9809 11887 9815 11913
rect 9841 11887 9847 11913
rect 12895 11881 12921 11887
rect 13231 11913 13257 11919
rect 13231 11881 13257 11887
rect 13287 11913 13313 11919
rect 13287 11881 13313 11887
rect 6791 11857 6817 11863
rect 6791 11825 6817 11831
rect 7687 11857 7713 11863
rect 7687 11825 7713 11831
rect 7799 11857 7825 11863
rect 10207 11857 10233 11863
rect 10711 11857 10737 11863
rect 8017 11831 8023 11857
rect 8049 11831 8055 11857
rect 9753 11831 9759 11857
rect 9785 11831 9791 11857
rect 10369 11831 10375 11857
rect 10401 11831 10407 11857
rect 7799 11825 7825 11831
rect 10207 11825 10233 11831
rect 10711 11825 10737 11831
rect 11047 11857 11073 11863
rect 11047 11825 11073 11831
rect 13007 11857 13033 11863
rect 13007 11825 13033 11831
rect 13399 11857 13425 11863
rect 14065 11831 14071 11857
rect 14097 11831 14103 11857
rect 13399 11825 13425 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 6231 11689 6257 11695
rect 6231 11657 6257 11663
rect 7183 11689 7209 11695
rect 7183 11657 7209 11663
rect 7295 11689 7321 11695
rect 11159 11689 11185 11695
rect 9809 11663 9815 11689
rect 9841 11663 9847 11689
rect 7295 11657 7321 11663
rect 11159 11657 11185 11663
rect 6903 11633 6929 11639
rect 6841 11607 6847 11633
rect 6873 11607 6879 11633
rect 6903 11601 6929 11607
rect 6959 11633 6985 11639
rect 6959 11601 6985 11607
rect 7071 11633 7097 11639
rect 7071 11601 7097 11607
rect 7351 11633 7377 11639
rect 10263 11633 10289 11639
rect 8409 11607 8415 11633
rect 8441 11607 8447 11633
rect 9025 11607 9031 11633
rect 9057 11607 9063 11633
rect 7351 11601 7377 11607
rect 10263 11601 10289 11607
rect 11103 11633 11129 11639
rect 11103 11601 11129 11607
rect 11215 11633 11241 11639
rect 11215 11601 11241 11607
rect 11439 11633 11465 11639
rect 11439 11601 11465 11607
rect 11495 11633 11521 11639
rect 11887 11633 11913 11639
rect 11713 11607 11719 11633
rect 11745 11607 11751 11633
rect 11495 11601 11521 11607
rect 11887 11601 11913 11607
rect 6287 11577 6313 11583
rect 6287 11545 6313 11551
rect 7015 11577 7041 11583
rect 10823 11577 10849 11583
rect 8297 11551 8303 11577
rect 8329 11551 8335 11577
rect 8969 11551 8975 11577
rect 9001 11551 9007 11577
rect 7015 11545 7041 11551
rect 10823 11545 10849 11551
rect 12111 11577 12137 11583
rect 12111 11545 12137 11551
rect 12223 11577 12249 11583
rect 12223 11545 12249 11551
rect 12391 11577 12417 11583
rect 12833 11551 12839 11577
rect 12865 11551 12871 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 12391 11545 12417 11551
rect 8807 11521 8833 11527
rect 8807 11489 8833 11495
rect 12279 11521 12305 11527
rect 14519 11521 14545 11527
rect 13225 11495 13231 11521
rect 13257 11495 13263 11521
rect 14289 11495 14295 11521
rect 14321 11495 14327 11521
rect 12279 11489 12305 11495
rect 14519 11489 14545 11495
rect 11439 11465 11465 11471
rect 11439 11433 11465 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 12111 11297 12137 11303
rect 12111 11265 12137 11271
rect 7071 11241 7097 11247
rect 11831 11241 11857 11247
rect 14631 11241 14657 11247
rect 11377 11215 11383 11241
rect 11409 11215 11415 11241
rect 13225 11215 13231 11241
rect 13257 11215 13263 11241
rect 14289 11215 14295 11241
rect 14321 11215 14327 11241
rect 7071 11209 7097 11215
rect 11831 11209 11857 11215
rect 14631 11209 14657 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 6959 11185 6985 11191
rect 6959 11153 6985 11159
rect 8135 11185 8161 11191
rect 8135 11153 8161 11159
rect 8359 11185 8385 11191
rect 8359 11153 8385 11159
rect 8415 11185 8441 11191
rect 8415 11153 8441 11159
rect 8807 11185 8833 11191
rect 8807 11153 8833 11159
rect 9647 11185 9673 11191
rect 9647 11153 9673 11159
rect 11159 11185 11185 11191
rect 11943 11185 11969 11191
rect 12391 11185 12417 11191
rect 11321 11159 11327 11185
rect 11353 11159 11359 11185
rect 12273 11159 12279 11185
rect 12305 11159 12311 11185
rect 11159 11153 11185 11159
rect 11943 11153 11969 11159
rect 12391 11153 12417 11159
rect 12503 11185 12529 11191
rect 12503 11153 12529 11159
rect 12889 11153 12895 11179
rect 12921 11153 12927 11179
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 6343 11129 6369 11135
rect 9031 11129 9057 11135
rect 6785 11103 6791 11129
rect 6817 11103 6823 11129
rect 10201 11103 10207 11129
rect 10233 11103 10239 11129
rect 10705 11103 10711 11129
rect 10737 11103 10743 11129
rect 6343 11097 6369 11103
rect 9031 11097 9057 11103
rect 6175 11073 6201 11079
rect 6175 11041 6201 11047
rect 8471 11073 8497 11079
rect 8471 11041 8497 11047
rect 9927 11073 9953 11079
rect 9927 11041 9953 11047
rect 10375 11073 10401 11079
rect 10375 11041 10401 11047
rect 10879 11073 10905 11079
rect 12335 11073 12361 11079
rect 11209 11047 11215 11073
rect 11241 11047 11247 11073
rect 10879 11041 10905 11047
rect 12335 11041 12361 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8079 10905 8105 10911
rect 12783 10905 12809 10911
rect 9193 10879 9199 10905
rect 9225 10879 9231 10905
rect 8079 10873 8105 10879
rect 12783 10873 12809 10879
rect 12839 10905 12865 10911
rect 12839 10873 12865 10879
rect 13175 10905 13201 10911
rect 13175 10873 13201 10879
rect 7855 10849 7881 10855
rect 12951 10849 12977 10855
rect 5889 10823 5895 10849
rect 5921 10823 5927 10849
rect 8913 10823 8919 10849
rect 8945 10823 8951 10849
rect 7855 10817 7881 10823
rect 12951 10817 12977 10823
rect 7183 10793 7209 10799
rect 5553 10767 5559 10793
rect 5585 10767 5591 10793
rect 7183 10761 7209 10767
rect 7575 10793 7601 10799
rect 7575 10761 7601 10767
rect 8247 10793 8273 10799
rect 12727 10793 12753 10799
rect 8353 10767 8359 10793
rect 8385 10767 8391 10793
rect 8689 10767 8695 10793
rect 8721 10767 8727 10793
rect 9137 10767 9143 10793
rect 9169 10767 9175 10793
rect 9585 10767 9591 10793
rect 9617 10767 9623 10793
rect 12609 10767 12615 10793
rect 12641 10767 12647 10793
rect 8247 10761 8273 10767
rect 12727 10761 12753 10767
rect 13119 10737 13145 10743
rect 6953 10711 6959 10737
rect 6985 10711 6991 10737
rect 11153 10711 11159 10737
rect 11185 10711 11191 10737
rect 13119 10705 13145 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7295 10457 7321 10463
rect 20007 10457 20033 10463
rect 7849 10431 7855 10457
rect 7881 10431 7887 10457
rect 13001 10431 13007 10457
rect 13033 10431 13039 10457
rect 7295 10425 7321 10431
rect 20007 10425 20033 10431
rect 6959 10401 6985 10407
rect 6959 10369 6985 10375
rect 7407 10401 7433 10407
rect 10655 10401 10681 10407
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 11153 10375 11159 10401
rect 11185 10375 11191 10401
rect 18937 10375 18943 10401
rect 18969 10375 18975 10401
rect 7407 10369 7433 10375
rect 10655 10369 10681 10375
rect 10879 10345 10905 10351
rect 10879 10313 10905 10319
rect 10991 10345 11017 10351
rect 10991 10313 11017 10319
rect 10823 10289 10849 10295
rect 7121 10263 7127 10289
rect 7153 10263 7159 10289
rect 7569 10263 7575 10289
rect 7601 10263 7607 10289
rect 10823 10257 10849 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 10207 10121 10233 10127
rect 10481 10095 10487 10121
rect 10513 10095 10519 10121
rect 10207 10089 10233 10095
rect 8695 10065 8721 10071
rect 7065 10039 7071 10065
rect 7097 10039 7103 10065
rect 10425 10039 10431 10065
rect 10457 10039 10463 10065
rect 12273 10039 12279 10065
rect 12305 10039 12311 10065
rect 8695 10033 8721 10039
rect 7239 10009 7265 10015
rect 7239 9977 7265 9983
rect 7407 10009 7433 10015
rect 7407 9977 7433 9983
rect 7911 10009 7937 10015
rect 7911 9977 7937 9983
rect 8191 10009 8217 10015
rect 8191 9977 8217 9983
rect 9367 10009 9393 10015
rect 9367 9977 9393 9983
rect 9479 10009 9505 10015
rect 11153 9983 11159 10009
rect 11185 9983 11191 10009
rect 11377 9983 11383 10009
rect 11409 9983 11415 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 9479 9977 9505 9983
rect 7625 9927 7631 9953
rect 7657 9927 7663 9953
rect 8857 9927 8863 9953
rect 8889 9927 8895 9953
rect 9977 9927 9983 9953
rect 10009 9927 10015 9953
rect 9535 9897 9561 9903
rect 9535 9865 9561 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 11495 9729 11521 9735
rect 11495 9697 11521 9703
rect 9423 9673 9449 9679
rect 11719 9673 11745 9679
rect 13847 9673 13873 9679
rect 8353 9647 8359 9673
rect 8385 9647 8391 9673
rect 9137 9647 9143 9673
rect 9169 9647 9175 9673
rect 9865 9647 9871 9673
rect 9897 9647 9903 9673
rect 12105 9647 12111 9673
rect 12137 9647 12143 9673
rect 9423 9641 9449 9647
rect 11719 9641 11745 9647
rect 13847 9641 13873 9647
rect 14071 9673 14097 9679
rect 14071 9641 14097 9647
rect 20007 9673 20033 9679
rect 20007 9641 20033 9647
rect 8807 9617 8833 9623
rect 8241 9591 8247 9617
rect 8273 9591 8279 9617
rect 8521 9591 8527 9617
rect 8553 9591 8559 9617
rect 8807 9585 8833 9591
rect 9255 9617 9281 9623
rect 11159 9617 11185 9623
rect 9753 9591 9759 9617
rect 9785 9591 9791 9617
rect 10313 9591 10319 9617
rect 10345 9591 10351 9617
rect 10705 9591 10711 9617
rect 10737 9591 10743 9617
rect 10929 9591 10935 9617
rect 10961 9591 10967 9617
rect 9255 9585 9281 9591
rect 11159 9585 11185 9591
rect 11327 9617 11353 9623
rect 11327 9585 11353 9591
rect 11383 9617 11409 9623
rect 11383 9585 11409 9591
rect 12447 9617 12473 9623
rect 12447 9585 12473 9591
rect 12615 9617 12641 9623
rect 12615 9585 12641 9591
rect 12727 9617 12753 9623
rect 12727 9585 12753 9591
rect 12951 9617 12977 9623
rect 12951 9585 12977 9591
rect 13063 9617 13089 9623
rect 14681 9591 14687 9617
rect 14713 9591 14719 9617
rect 15017 9591 15023 9617
rect 15049 9591 15055 9617
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 13063 9585 13089 9591
rect 13623 9561 13649 9567
rect 9865 9535 9871 9561
rect 9897 9535 9903 9561
rect 12273 9535 12279 9561
rect 12305 9535 12311 9561
rect 13623 9529 13649 9535
rect 13735 9561 13761 9567
rect 13735 9529 13761 9535
rect 13903 9561 13929 9567
rect 14793 9535 14799 9561
rect 14825 9535 14831 9561
rect 13903 9529 13929 9535
rect 8695 9505 8721 9511
rect 8695 9473 8721 9479
rect 8751 9505 8777 9511
rect 8751 9473 8777 9479
rect 12559 9505 12585 9511
rect 12559 9473 12585 9479
rect 13007 9505 13033 9511
rect 13007 9473 13033 9479
rect 13175 9505 13201 9511
rect 13175 9473 13201 9479
rect 13455 9505 13481 9511
rect 13455 9473 13481 9479
rect 14127 9505 14153 9511
rect 14127 9473 14153 9479
rect 14183 9505 14209 9511
rect 15129 9479 15135 9505
rect 15161 9479 15167 9505
rect 14183 9473 14209 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 13007 9337 13033 9343
rect 9249 9311 9255 9337
rect 9281 9311 9287 9337
rect 11265 9311 11271 9337
rect 11297 9311 11303 9337
rect 13007 9305 13033 9311
rect 10487 9281 10513 9287
rect 10487 9249 10513 9255
rect 11495 9281 11521 9287
rect 11495 9249 11521 9255
rect 12167 9281 12193 9287
rect 12167 9249 12193 9255
rect 12279 9281 12305 9287
rect 12279 9249 12305 9255
rect 12671 9281 12697 9287
rect 12671 9249 12697 9255
rect 12727 9281 12753 9287
rect 12727 9249 12753 9255
rect 12951 9281 12977 9287
rect 13785 9255 13791 9281
rect 13817 9255 13823 9281
rect 12951 9249 12977 9255
rect 7407 9225 7433 9231
rect 5721 9199 5727 9225
rect 5753 9199 5759 9225
rect 6113 9199 6119 9225
rect 6145 9199 6151 9225
rect 7407 9193 7433 9199
rect 8695 9225 8721 9231
rect 8695 9193 8721 9199
rect 8975 9225 9001 9231
rect 8975 9193 9001 9199
rect 9423 9225 9449 9231
rect 10935 9225 10961 9231
rect 10761 9199 10767 9225
rect 10793 9199 10799 9225
rect 9423 9193 9449 9199
rect 10935 9193 10961 9199
rect 11999 9225 12025 9231
rect 11999 9193 12025 9199
rect 12055 9225 12081 9231
rect 12055 9193 12081 9199
rect 12559 9225 12585 9231
rect 12559 9193 12585 9199
rect 13119 9225 13145 9231
rect 13393 9199 13399 9225
rect 13425 9199 13431 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 13119 9193 13145 9199
rect 12111 9169 12137 9175
rect 7177 9143 7183 9169
rect 7209 9143 7215 9169
rect 14849 9143 14855 9169
rect 14881 9143 14887 9169
rect 12111 9137 12137 9143
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 8583 8945 8609 8951
rect 8583 8913 8609 8919
rect 9423 8945 9449 8951
rect 9423 8913 9449 8919
rect 11495 8945 11521 8951
rect 11495 8913 11521 8919
rect 967 8889 993 8895
rect 967 8857 993 8863
rect 8471 8889 8497 8895
rect 10207 8889 10233 8895
rect 9249 8863 9255 8889
rect 9281 8863 9287 8889
rect 9585 8863 9591 8889
rect 9617 8863 9623 8889
rect 8471 8857 8497 8863
rect 10207 8857 10233 8863
rect 10655 8889 10681 8895
rect 10655 8857 10681 8863
rect 11439 8889 11465 8895
rect 20007 8889 20033 8895
rect 12049 8863 12055 8889
rect 12081 8863 12087 8889
rect 13113 8863 13119 8889
rect 13145 8863 13151 8889
rect 11439 8857 11465 8863
rect 20007 8857 20033 8863
rect 7295 8833 7321 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 7295 8801 7321 8807
rect 7687 8833 7713 8839
rect 7687 8801 7713 8807
rect 7855 8833 7881 8839
rect 9087 8833 9113 8839
rect 9927 8833 9953 8839
rect 7961 8807 7967 8833
rect 7993 8807 7999 8833
rect 9697 8807 9703 8833
rect 9729 8807 9735 8833
rect 7855 8801 7881 8807
rect 9087 8801 9113 8807
rect 9927 8801 9953 8807
rect 10711 8833 10737 8839
rect 10711 8801 10737 8807
rect 10823 8833 10849 8839
rect 10823 8801 10849 8807
rect 11103 8833 11129 8839
rect 13231 8833 13257 8839
rect 11321 8807 11327 8833
rect 11353 8807 11359 8833
rect 11713 8807 11719 8833
rect 11745 8807 11751 8833
rect 11103 8801 11129 8807
rect 13231 8801 13257 8807
rect 13511 8833 13537 8839
rect 13511 8801 13537 8807
rect 13735 8833 13761 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 13735 8801 13761 8807
rect 7351 8777 7377 8783
rect 9311 8777 9337 8783
rect 8913 8751 8919 8777
rect 8945 8751 8951 8777
rect 7351 8745 7377 8751
rect 9311 8745 9337 8751
rect 11047 8777 11073 8783
rect 11047 8745 11073 8751
rect 13455 8777 13481 8783
rect 13455 8745 13481 8751
rect 13791 8777 13817 8783
rect 13791 8745 13817 8751
rect 13903 8777 13929 8783
rect 13903 8745 13929 8751
rect 7463 8721 7489 8727
rect 7463 8689 7489 8695
rect 7743 8721 7769 8727
rect 7743 8689 7769 8695
rect 7799 8721 7825 8727
rect 10935 8721 10961 8727
rect 8745 8695 8751 8721
rect 8777 8695 8783 8721
rect 7799 8689 7825 8695
rect 10935 8689 10961 8695
rect 13343 8721 13369 8727
rect 13343 8689 13369 8695
rect 14071 8721 14097 8727
rect 14071 8689 14097 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7967 8553 7993 8559
rect 7967 8521 7993 8527
rect 8247 8553 8273 8559
rect 8247 8521 8273 8527
rect 10655 8553 10681 8559
rect 10655 8521 10681 8527
rect 12839 8553 12865 8559
rect 12839 8521 12865 8527
rect 7351 8497 7377 8503
rect 6785 8471 6791 8497
rect 6817 8471 6823 8497
rect 7351 8465 7377 8471
rect 7407 8497 7433 8503
rect 9249 8471 9255 8497
rect 9281 8471 9287 8497
rect 13393 8471 13399 8497
rect 13425 8471 13431 8497
rect 7407 8465 7433 8471
rect 7519 8441 7545 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7177 8415 7183 8441
rect 7209 8415 7215 8441
rect 7519 8409 7545 8415
rect 7743 8441 7769 8447
rect 7743 8409 7769 8415
rect 7799 8441 7825 8447
rect 7799 8409 7825 8415
rect 7911 8441 7937 8447
rect 9137 8415 9143 8441
rect 9169 8415 9175 8441
rect 13001 8415 13007 8441
rect 13033 8415 13039 8441
rect 7911 8409 7937 8415
rect 7855 8385 7881 8391
rect 5721 8359 5727 8385
rect 5753 8359 5759 8385
rect 7855 8353 7881 8359
rect 10711 8385 10737 8391
rect 10711 8353 10737 8359
rect 10767 8385 10793 8391
rect 14457 8359 14463 8385
rect 14489 8359 14495 8385
rect 10767 8353 10793 8359
rect 967 8329 993 8335
rect 967 8297 993 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 11551 8161 11577 8167
rect 11551 8129 11577 8135
rect 13567 8161 13593 8167
rect 13567 8129 13593 8135
rect 11663 8105 11689 8111
rect 1017 8079 1023 8105
rect 1049 8079 1055 8105
rect 11663 8073 11689 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 7239 8049 7265 8055
rect 2137 8023 2143 8049
rect 2169 8023 2175 8049
rect 7239 8017 7265 8023
rect 7687 8049 7713 8055
rect 7687 8017 7713 8023
rect 7799 8049 7825 8055
rect 13729 8023 13735 8049
rect 13761 8023 13767 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 7799 8017 7825 8023
rect 7407 7993 7433 7999
rect 7407 7961 7433 7967
rect 7519 7993 7545 7999
rect 7519 7961 7545 7967
rect 7295 7937 7321 7943
rect 7295 7905 7321 7911
rect 7575 7937 7601 7943
rect 7575 7905 7601 7911
rect 8919 7937 8945 7943
rect 13623 7937 13649 7943
rect 11377 7911 11383 7937
rect 11409 7911 11415 7937
rect 8919 7905 8945 7911
rect 13623 7905 13649 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 14519 7769 14545 7775
rect 14519 7737 14545 7743
rect 8807 7713 8833 7719
rect 6897 7687 6903 7713
rect 6929 7687 6935 7713
rect 9137 7687 9143 7713
rect 9169 7687 9175 7713
rect 10985 7687 10991 7713
rect 11017 7687 11023 7713
rect 8807 7681 8833 7687
rect 7519 7657 7545 7663
rect 7233 7631 7239 7657
rect 7265 7631 7271 7657
rect 7519 7625 7545 7631
rect 8919 7657 8945 7663
rect 9249 7631 9255 7657
rect 9281 7631 9287 7657
rect 11377 7631 11383 7657
rect 11409 7631 11415 7657
rect 12833 7631 12839 7657
rect 12865 7631 12871 7657
rect 8919 7625 8945 7631
rect 8863 7601 8889 7607
rect 11607 7601 11633 7607
rect 5833 7575 5839 7601
rect 5865 7575 5871 7601
rect 9921 7575 9927 7601
rect 9953 7575 9959 7601
rect 13225 7575 13231 7601
rect 13257 7575 13263 7601
rect 14289 7575 14295 7601
rect 14321 7575 14327 7601
rect 8863 7569 8889 7575
rect 11607 7569 11633 7575
rect 9031 7545 9057 7551
rect 9031 7513 9057 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9031 7377 9057 7383
rect 9031 7345 9057 7351
rect 9983 7377 10009 7383
rect 9983 7345 10009 7351
rect 10879 7377 10905 7383
rect 10879 7345 10905 7351
rect 11439 7377 11465 7383
rect 11439 7345 11465 7351
rect 11719 7377 11745 7383
rect 11719 7345 11745 7351
rect 13343 7377 13369 7383
rect 13343 7345 13369 7351
rect 9367 7321 9393 7327
rect 7737 7295 7743 7321
rect 7769 7295 7775 7321
rect 8801 7295 8807 7321
rect 8833 7295 8839 7321
rect 9193 7295 9199 7321
rect 9225 7295 9231 7321
rect 9367 7289 9393 7295
rect 9591 7321 9617 7327
rect 11383 7321 11409 7327
rect 10145 7295 10151 7321
rect 10177 7295 10183 7321
rect 11041 7295 11047 7321
rect 11073 7295 11079 7321
rect 13225 7295 13231 7321
rect 13257 7295 13263 7321
rect 9591 7289 9617 7295
rect 11383 7289 11409 7295
rect 9759 7265 9785 7271
rect 7401 7239 7407 7265
rect 7433 7239 7439 7265
rect 9759 7233 9785 7239
rect 11271 7265 11297 7271
rect 11271 7233 11297 7239
rect 11831 7265 11857 7271
rect 11937 7239 11943 7265
rect 11969 7239 11975 7265
rect 13169 7239 13175 7265
rect 13201 7239 13207 7265
rect 11831 7233 11857 7239
rect 8975 7209 9001 7215
rect 8975 7177 9001 7183
rect 9255 7209 9281 7215
rect 9255 7177 9281 7183
rect 9535 7209 9561 7215
rect 9535 7177 9561 7183
rect 9703 7209 9729 7215
rect 9703 7177 9729 7183
rect 11215 7209 11241 7215
rect 11215 7177 11241 7183
rect 11663 7209 11689 7215
rect 11663 7177 11689 7183
rect 10095 7153 10121 7159
rect 10095 7121 10121 7127
rect 10375 7153 10401 7159
rect 10375 7121 10401 7127
rect 10991 7153 11017 7159
rect 10991 7121 11017 7127
rect 12391 7153 12417 7159
rect 12391 7121 12417 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 7575 6985 7601 6991
rect 7575 6953 7601 6959
rect 12671 6985 12697 6991
rect 12671 6953 12697 6959
rect 12615 6929 12641 6935
rect 6953 6903 6959 6929
rect 6985 6903 6991 6929
rect 9081 6903 9087 6929
rect 9113 6903 9119 6929
rect 11209 6903 11215 6929
rect 11241 6903 11247 6929
rect 12615 6897 12641 6903
rect 10431 6873 10457 6879
rect 7345 6847 7351 6873
rect 7377 6847 7383 6873
rect 8745 6847 8751 6873
rect 8777 6847 8783 6873
rect 10313 6847 10319 6873
rect 10345 6847 10351 6873
rect 10431 6841 10457 6847
rect 10543 6873 10569 6879
rect 10873 6847 10879 6873
rect 10905 6847 10911 6873
rect 12777 6847 12783 6873
rect 12809 6847 12815 6873
rect 10543 6841 10569 6847
rect 5889 6791 5895 6817
rect 5921 6791 5927 6817
rect 10145 6791 10151 6817
rect 10177 6791 10183 6817
rect 12273 6791 12279 6817
rect 12305 6791 12311 6817
rect 10599 6761 10625 6767
rect 10599 6729 10625 6735
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 8807 6537 8833 6543
rect 13119 6537 13145 6543
rect 9305 6511 9311 6537
rect 9337 6511 9343 6537
rect 10369 6511 10375 6537
rect 10401 6511 10407 6537
rect 11769 6511 11775 6537
rect 11801 6511 11807 6537
rect 12833 6511 12839 6537
rect 12865 6511 12871 6537
rect 8807 6505 8833 6511
rect 13119 6505 13145 6511
rect 8913 6455 8919 6481
rect 8945 6455 8951 6481
rect 11433 6455 11439 6481
rect 11465 6455 11471 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8969 2143 8975 2169
rect 9001 2143 9007 2169
rect 10369 2143 10375 2169
rect 10401 2143 10407 2169
rect 12833 2143 12839 2169
rect 12865 2143 12871 2169
rect 9255 2057 9281 2063
rect 9255 2025 9281 2031
rect 10711 2057 10737 2063
rect 10711 2025 10737 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 9865 1751 9871 1777
rect 9897 1751 9903 1777
rect 10817 1751 10823 1777
rect 10849 1751 10855 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 9591 1665 9617 1671
rect 9591 1633 9617 1639
rect 11215 1665 11241 1671
rect 11215 1633 11241 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 11047 19111 11073 19137
rect 12783 19111 12809 19137
rect 8807 18999 8833 19025
rect 10543 18999 10569 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9199 18719 9225 18745
rect 10151 18719 10177 18745
rect 13399 18719 13425 18745
rect 8807 18607 8833 18633
rect 12895 18607 12921 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 20119 17319 20145 17345
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 8527 14351 8553 14377
rect 12111 14351 12137 14377
rect 7127 14295 7153 14321
rect 10711 14295 10737 14321
rect 11047 14295 11073 14321
rect 12335 14295 12361 14321
rect 7463 14239 7489 14265
rect 8863 14183 8889 14209
rect 9087 14183 9113 14209
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8191 14015 8217 14041
rect 10879 14015 10905 14041
rect 8751 13959 8777 13985
rect 10711 13959 10737 13985
rect 11271 13959 11297 13985
rect 8135 13903 8161 13929
rect 8247 13903 8273 13929
rect 8471 13903 8497 13929
rect 8695 13903 8721 13929
rect 9031 13903 9057 13929
rect 10823 13903 10849 13929
rect 10935 13903 10961 13929
rect 11215 13903 11241 13929
rect 9423 13847 9449 13873
rect 10487 13847 10513 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 8527 13567 8553 13593
rect 9199 13567 9225 13593
rect 9535 13567 9561 13593
rect 12895 13567 12921 13593
rect 7127 13511 7153 13537
rect 8807 13511 8833 13537
rect 8919 13511 8945 13537
rect 9479 13511 9505 13537
rect 9591 13511 9617 13537
rect 9815 13511 9841 13537
rect 10095 13511 10121 13537
rect 10375 13511 10401 13537
rect 11439 13511 11465 13537
rect 7463 13455 7489 13481
rect 8695 13455 8721 13481
rect 8751 13455 8777 13481
rect 10151 13455 10177 13481
rect 11831 13455 11857 13481
rect 9703 13399 9729 13425
rect 10039 13399 10065 13425
rect 13119 13399 13145 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8863 13231 8889 13257
rect 10879 13231 10905 13257
rect 11607 13231 11633 13257
rect 8695 13175 8721 13201
rect 12671 13175 12697 13201
rect 8807 13119 8833 13145
rect 8919 13119 8945 13145
rect 8975 13119 9001 13145
rect 11047 13119 11073 13145
rect 11551 13119 11577 13145
rect 11663 13119 11689 13145
rect 12615 13119 12641 13145
rect 11439 13063 11465 13089
rect 11215 13007 11241 13033
rect 11327 13007 11353 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 8135 12839 8161 12865
rect 9927 12839 9953 12865
rect 10711 12839 10737 12865
rect 9031 12783 9057 12809
rect 12447 12783 12473 12809
rect 12671 12783 12697 12809
rect 8191 12727 8217 12753
rect 10991 12727 11017 12753
rect 8919 12671 8945 12697
rect 9871 12671 9897 12697
rect 10655 12671 10681 12697
rect 11383 12671 11409 12697
rect 7911 12615 7937 12641
rect 8135 12615 8161 12641
rect 8359 12615 8385 12641
rect 8527 12615 8553 12641
rect 8975 12615 9001 12641
rect 9927 12615 9953 12641
rect 10711 12615 10737 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8863 12447 8889 12473
rect 11663 12447 11689 12473
rect 12111 12447 12137 12473
rect 8247 12391 8273 12417
rect 8919 12391 8945 12417
rect 10263 12391 10289 12417
rect 6455 12335 6481 12361
rect 8359 12335 8385 12361
rect 9647 12335 9673 12361
rect 10151 12335 10177 12361
rect 6847 12279 6873 12305
rect 7911 12279 7937 12305
rect 9423 12279 9449 12305
rect 11383 12279 11409 12305
rect 11887 12279 11913 12305
rect 8807 12223 8833 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 967 11999 993 12025
rect 4999 11999 5025 12025
rect 8191 11999 8217 12025
rect 8415 11999 8441 12025
rect 9591 11999 9617 12025
rect 10655 11999 10681 12025
rect 13063 11999 13089 12025
rect 20007 11999 20033 12025
rect 2143 11943 2169 11969
rect 6399 11943 6425 11969
rect 7855 11943 7881 11969
rect 8303 11943 8329 11969
rect 8527 11943 8553 11969
rect 9367 11943 9393 11969
rect 9983 11943 10009 11969
rect 11047 11943 11073 11969
rect 13959 11943 13985 11969
rect 18831 11943 18857 11969
rect 6063 11887 6089 11913
rect 8583 11887 8609 11913
rect 8975 11887 9001 11913
rect 9815 11887 9841 11913
rect 12895 11887 12921 11913
rect 13231 11887 13257 11913
rect 13287 11887 13313 11913
rect 6791 11831 6817 11857
rect 7687 11831 7713 11857
rect 7799 11831 7825 11857
rect 8023 11831 8049 11857
rect 9759 11831 9785 11857
rect 10207 11831 10233 11857
rect 10375 11831 10401 11857
rect 10711 11831 10737 11857
rect 11047 11831 11073 11857
rect 13007 11831 13033 11857
rect 13399 11831 13425 11857
rect 14071 11831 14097 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 6231 11663 6257 11689
rect 7183 11663 7209 11689
rect 7295 11663 7321 11689
rect 9815 11663 9841 11689
rect 11159 11663 11185 11689
rect 6847 11607 6873 11633
rect 6903 11607 6929 11633
rect 6959 11607 6985 11633
rect 7071 11607 7097 11633
rect 7351 11607 7377 11633
rect 8415 11607 8441 11633
rect 9031 11607 9057 11633
rect 10263 11607 10289 11633
rect 11103 11607 11129 11633
rect 11215 11607 11241 11633
rect 11439 11607 11465 11633
rect 11495 11607 11521 11633
rect 11719 11607 11745 11633
rect 11887 11607 11913 11633
rect 6287 11551 6313 11577
rect 7015 11551 7041 11577
rect 8303 11551 8329 11577
rect 8975 11551 9001 11577
rect 10823 11551 10849 11577
rect 12111 11551 12137 11577
rect 12223 11551 12249 11577
rect 12391 11551 12417 11577
rect 12839 11551 12865 11577
rect 18831 11551 18857 11577
rect 8807 11495 8833 11521
rect 12279 11495 12305 11521
rect 13231 11495 13257 11521
rect 14295 11495 14321 11521
rect 14519 11495 14545 11521
rect 11439 11439 11465 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 12111 11271 12137 11297
rect 7071 11215 7097 11241
rect 11383 11215 11409 11241
rect 11831 11215 11857 11241
rect 13231 11215 13257 11241
rect 14295 11215 14321 11241
rect 14631 11215 14657 11241
rect 20007 11215 20033 11241
rect 6959 11159 6985 11185
rect 8135 11159 8161 11185
rect 8359 11159 8385 11185
rect 8415 11159 8441 11185
rect 8807 11159 8833 11185
rect 9647 11159 9673 11185
rect 11159 11159 11185 11185
rect 11327 11159 11353 11185
rect 11943 11159 11969 11185
rect 12279 11159 12305 11185
rect 12391 11159 12417 11185
rect 12503 11159 12529 11185
rect 12895 11153 12921 11179
rect 18831 11159 18857 11185
rect 6343 11103 6369 11129
rect 6791 11103 6817 11129
rect 9031 11103 9057 11129
rect 10207 11103 10233 11129
rect 10711 11103 10737 11129
rect 6175 11047 6201 11073
rect 8471 11047 8497 11073
rect 9927 11047 9953 11073
rect 10375 11047 10401 11073
rect 10879 11047 10905 11073
rect 11215 11047 11241 11073
rect 12335 11047 12361 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8079 10879 8105 10905
rect 9199 10879 9225 10905
rect 12783 10879 12809 10905
rect 12839 10879 12865 10905
rect 13175 10879 13201 10905
rect 5895 10823 5921 10849
rect 7855 10823 7881 10849
rect 8919 10823 8945 10849
rect 12951 10823 12977 10849
rect 5559 10767 5585 10793
rect 7183 10767 7209 10793
rect 7575 10767 7601 10793
rect 8247 10767 8273 10793
rect 8359 10767 8385 10793
rect 8695 10767 8721 10793
rect 9143 10767 9169 10793
rect 9591 10767 9617 10793
rect 12615 10767 12641 10793
rect 12727 10767 12753 10793
rect 6959 10711 6985 10737
rect 11159 10711 11185 10737
rect 13119 10711 13145 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7295 10431 7321 10457
rect 7855 10431 7881 10457
rect 13007 10431 13033 10457
rect 20007 10431 20033 10457
rect 6959 10375 6985 10401
rect 7407 10375 7433 10401
rect 10039 10375 10065 10401
rect 10655 10375 10681 10401
rect 11159 10375 11185 10401
rect 18943 10375 18969 10401
rect 10879 10319 10905 10345
rect 10991 10319 11017 10345
rect 7127 10263 7153 10289
rect 7575 10263 7601 10289
rect 10823 10263 10849 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 10207 10095 10233 10121
rect 10487 10095 10513 10121
rect 7071 10039 7097 10065
rect 8695 10039 8721 10065
rect 10431 10039 10457 10065
rect 12279 10039 12305 10065
rect 7239 9983 7265 10009
rect 7407 9983 7433 10009
rect 7911 9983 7937 10009
rect 8191 9983 8217 10009
rect 9367 9983 9393 10009
rect 9479 9983 9505 10009
rect 11159 9983 11185 10009
rect 11383 9983 11409 10009
rect 18831 9983 18857 10009
rect 7631 9927 7657 9953
rect 8863 9927 8889 9953
rect 9983 9927 10009 9953
rect 9535 9871 9561 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 11495 9703 11521 9729
rect 8359 9647 8385 9673
rect 9143 9647 9169 9673
rect 9423 9647 9449 9673
rect 9871 9647 9897 9673
rect 11719 9647 11745 9673
rect 12111 9647 12137 9673
rect 13847 9647 13873 9673
rect 14071 9647 14097 9673
rect 20007 9647 20033 9673
rect 8247 9591 8273 9617
rect 8527 9591 8553 9617
rect 8807 9591 8833 9617
rect 9255 9591 9281 9617
rect 9759 9591 9785 9617
rect 10319 9591 10345 9617
rect 10711 9591 10737 9617
rect 10935 9591 10961 9617
rect 11159 9591 11185 9617
rect 11327 9591 11353 9617
rect 11383 9591 11409 9617
rect 12447 9591 12473 9617
rect 12615 9591 12641 9617
rect 12727 9591 12753 9617
rect 12951 9591 12977 9617
rect 13063 9591 13089 9617
rect 14687 9591 14713 9617
rect 15023 9591 15049 9617
rect 18831 9591 18857 9617
rect 9871 9535 9897 9561
rect 12279 9535 12305 9561
rect 13623 9535 13649 9561
rect 13735 9535 13761 9561
rect 13903 9535 13929 9561
rect 14799 9535 14825 9561
rect 8695 9479 8721 9505
rect 8751 9479 8777 9505
rect 12559 9479 12585 9505
rect 13007 9479 13033 9505
rect 13175 9479 13201 9505
rect 13455 9479 13481 9505
rect 14127 9479 14153 9505
rect 14183 9479 14209 9505
rect 15135 9479 15161 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 9255 9311 9281 9337
rect 11271 9311 11297 9337
rect 13007 9311 13033 9337
rect 10487 9255 10513 9281
rect 11495 9255 11521 9281
rect 12167 9255 12193 9281
rect 12279 9255 12305 9281
rect 12671 9255 12697 9281
rect 12727 9255 12753 9281
rect 12951 9255 12977 9281
rect 13791 9255 13817 9281
rect 5727 9199 5753 9225
rect 6119 9199 6145 9225
rect 7407 9199 7433 9225
rect 8695 9199 8721 9225
rect 8975 9199 9001 9225
rect 9423 9199 9449 9225
rect 10767 9199 10793 9225
rect 10935 9199 10961 9225
rect 11999 9199 12025 9225
rect 12055 9199 12081 9225
rect 12559 9199 12585 9225
rect 13119 9199 13145 9225
rect 13399 9199 13425 9225
rect 18831 9199 18857 9225
rect 7183 9143 7209 9169
rect 12111 9143 12137 9169
rect 14855 9143 14881 9169
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 8583 8919 8609 8945
rect 9423 8919 9449 8945
rect 11495 8919 11521 8945
rect 967 8863 993 8889
rect 8471 8863 8497 8889
rect 9255 8863 9281 8889
rect 9591 8863 9617 8889
rect 10207 8863 10233 8889
rect 10655 8863 10681 8889
rect 11439 8863 11465 8889
rect 12055 8863 12081 8889
rect 13119 8863 13145 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 7295 8807 7321 8833
rect 7687 8807 7713 8833
rect 7855 8807 7881 8833
rect 7967 8807 7993 8833
rect 9087 8807 9113 8833
rect 9703 8807 9729 8833
rect 9927 8807 9953 8833
rect 10711 8807 10737 8833
rect 10823 8807 10849 8833
rect 11103 8807 11129 8833
rect 11327 8807 11353 8833
rect 11719 8807 11745 8833
rect 13231 8807 13257 8833
rect 13511 8807 13537 8833
rect 13735 8807 13761 8833
rect 18831 8807 18857 8833
rect 7351 8751 7377 8777
rect 8919 8751 8945 8777
rect 9311 8751 9337 8777
rect 11047 8751 11073 8777
rect 13455 8751 13481 8777
rect 13791 8751 13817 8777
rect 13903 8751 13929 8777
rect 7463 8695 7489 8721
rect 7743 8695 7769 8721
rect 7799 8695 7825 8721
rect 8751 8695 8777 8721
rect 10935 8695 10961 8721
rect 13343 8695 13369 8721
rect 14071 8695 14097 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7967 8527 7993 8553
rect 8247 8527 8273 8553
rect 10655 8527 10681 8553
rect 12839 8527 12865 8553
rect 6791 8471 6817 8497
rect 7351 8471 7377 8497
rect 7407 8471 7433 8497
rect 9255 8471 9281 8497
rect 13399 8471 13425 8497
rect 2143 8415 2169 8441
rect 7183 8415 7209 8441
rect 7519 8415 7545 8441
rect 7743 8415 7769 8441
rect 7799 8415 7825 8441
rect 7911 8415 7937 8441
rect 9143 8415 9169 8441
rect 13007 8415 13033 8441
rect 5727 8359 5753 8385
rect 7855 8359 7881 8385
rect 10711 8359 10737 8385
rect 10767 8359 10793 8385
rect 14463 8359 14489 8385
rect 967 8303 993 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 11551 8135 11577 8161
rect 13567 8135 13593 8161
rect 1023 8079 1049 8105
rect 11663 8079 11689 8105
rect 20007 8079 20033 8105
rect 2143 8023 2169 8049
rect 7239 8023 7265 8049
rect 7687 8023 7713 8049
rect 7799 8023 7825 8049
rect 13735 8023 13761 8049
rect 18831 8023 18857 8049
rect 7407 7967 7433 7993
rect 7519 7967 7545 7993
rect 7295 7911 7321 7937
rect 7575 7911 7601 7937
rect 8919 7911 8945 7937
rect 11383 7911 11409 7937
rect 13623 7911 13649 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 14519 7743 14545 7769
rect 6903 7687 6929 7713
rect 8807 7687 8833 7713
rect 9143 7687 9169 7713
rect 10991 7687 11017 7713
rect 7239 7631 7265 7657
rect 7519 7631 7545 7657
rect 8919 7631 8945 7657
rect 9255 7631 9281 7657
rect 11383 7631 11409 7657
rect 12839 7631 12865 7657
rect 5839 7575 5865 7601
rect 8863 7575 8889 7601
rect 9927 7575 9953 7601
rect 11607 7575 11633 7601
rect 13231 7575 13257 7601
rect 14295 7575 14321 7601
rect 9031 7519 9057 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9031 7351 9057 7377
rect 9983 7351 10009 7377
rect 10879 7351 10905 7377
rect 11439 7351 11465 7377
rect 11719 7351 11745 7377
rect 13343 7351 13369 7377
rect 7743 7295 7769 7321
rect 8807 7295 8833 7321
rect 9199 7295 9225 7321
rect 9367 7295 9393 7321
rect 9591 7295 9617 7321
rect 10151 7295 10177 7321
rect 11047 7295 11073 7321
rect 11383 7295 11409 7321
rect 13231 7295 13257 7321
rect 7407 7239 7433 7265
rect 9759 7239 9785 7265
rect 11271 7239 11297 7265
rect 11831 7239 11857 7265
rect 11943 7239 11969 7265
rect 13175 7239 13201 7265
rect 8975 7183 9001 7209
rect 9255 7183 9281 7209
rect 9535 7183 9561 7209
rect 9703 7183 9729 7209
rect 11215 7183 11241 7209
rect 11663 7183 11689 7209
rect 10095 7127 10121 7153
rect 10375 7127 10401 7153
rect 10991 7127 11017 7153
rect 12391 7127 12417 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 7575 6959 7601 6985
rect 12671 6959 12697 6985
rect 6959 6903 6985 6929
rect 9087 6903 9113 6929
rect 11215 6903 11241 6929
rect 12615 6903 12641 6929
rect 7351 6847 7377 6873
rect 8751 6847 8777 6873
rect 10319 6847 10345 6873
rect 10431 6847 10457 6873
rect 10543 6847 10569 6873
rect 10879 6847 10905 6873
rect 12783 6847 12809 6873
rect 5895 6791 5921 6817
rect 10151 6791 10177 6817
rect 12279 6791 12305 6817
rect 10599 6735 10625 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8807 6511 8833 6537
rect 9311 6511 9337 6537
rect 10375 6511 10401 6537
rect 11775 6511 11801 6537
rect 12839 6511 12865 6537
rect 13119 6511 13145 6537
rect 8919 6455 8945 6481
rect 11439 6455 11465 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8975 2143 9001 2169
rect 10375 2143 10401 2169
rect 12839 2143 12865 2169
rect 9255 2031 9281 2057
rect 10711 2031 10737 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 12783 1807 12809 1833
rect 9871 1751 9897 1777
rect 10823 1751 10849 1777
rect 12279 1751 12305 1777
rect 9591 1639 9617 1665
rect 11215 1639 11241 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 8736 20600 8792 21000
rect 9744 20600 9800 21000
rect 10416 20600 10472 21000
rect 11424 20600 11480 21000
rect 12768 20600 12824 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8414 18746 8442 20600
rect 8750 19138 8778 20600
rect 9758 19306 9786 20600
rect 9758 19278 10178 19306
rect 8750 19105 8778 19110
rect 9310 19138 9338 19143
rect 9310 19091 9338 19110
rect 8806 19026 8834 19031
rect 8414 18713 8442 18718
rect 8526 19025 8834 19026
rect 8526 18999 8807 19025
rect 8833 18999 8834 19025
rect 8526 18998 8834 18999
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 8526 14378 8554 18998
rect 8806 18993 8834 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9198 18746 9226 18751
rect 9198 18699 9226 18718
rect 10150 18745 10178 19278
rect 10430 19138 10458 20600
rect 10430 19105 10458 19110
rect 11046 19138 11074 19143
rect 11046 19091 11074 19110
rect 11438 19138 11466 20600
rect 12782 19306 12810 20600
rect 12782 19273 12810 19278
rect 13398 19306 13426 19311
rect 11438 19105 11466 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 10150 18719 10151 18745
rect 10177 18719 10178 18745
rect 10150 18713 10178 18719
rect 10542 19025 10570 19031
rect 10542 18999 10543 19025
rect 10569 18999 10570 19025
rect 8806 18633 8834 18639
rect 8806 18607 8807 18633
rect 8833 18607 8834 18633
rect 8526 14377 8778 14378
rect 8526 14351 8527 14377
rect 8553 14351 8778 14377
rect 8526 14350 8778 14351
rect 8526 14345 8554 14350
rect 7126 14321 7154 14327
rect 7126 14295 7127 14321
rect 7153 14295 7154 14321
rect 7126 14210 7154 14295
rect 7462 14266 7490 14271
rect 7462 14219 7490 14238
rect 8190 14266 8218 14271
rect 2086 14154 2114 14159
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 2086 11522 2114 14126
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 7126 13537 7154 14182
rect 8190 14041 8218 14238
rect 8190 14015 8191 14041
rect 8217 14015 8218 14041
rect 8190 14009 8218 14015
rect 8750 13985 8778 14350
rect 8750 13959 8751 13985
rect 8777 13959 8778 13985
rect 8750 13953 8778 13959
rect 8134 13929 8162 13935
rect 8134 13903 8135 13929
rect 8161 13903 8162 13929
rect 8134 13594 8162 13903
rect 8246 13930 8274 13935
rect 8246 13883 8274 13902
rect 8470 13929 8498 13935
rect 8470 13903 8471 13929
rect 8497 13903 8498 13929
rect 8134 13561 8162 13566
rect 7126 13511 7127 13537
rect 7153 13511 7154 13537
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6454 12418 6482 12423
rect 6454 12362 6482 12390
rect 7126 12418 7154 13511
rect 7462 13482 7490 13487
rect 8470 13454 8498 13903
rect 8694 13930 8722 13935
rect 8694 13883 8722 13902
rect 8806 13818 8834 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 10542 15974 10570 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 13398 18745 13426 19278
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 13398 18719 13399 18745
rect 13425 18719 13426 18745
rect 13398 18713 13426 18719
rect 10486 15946 10570 15974
rect 12110 15946 12306 15974
rect 12894 18633 12922 18639
rect 12894 18607 12895 18633
rect 12921 18607 12922 18633
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 8862 14210 8890 14215
rect 9086 14210 9114 14215
rect 8890 14209 9114 14210
rect 8890 14183 9087 14209
rect 9113 14183 9114 14209
rect 8890 14182 9114 14183
rect 8862 14163 8890 14182
rect 9030 13930 9058 14182
rect 9086 14177 9114 14182
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9030 13929 9226 13930
rect 9030 13903 9031 13929
rect 9057 13903 9226 13929
rect 9030 13902 9226 13903
rect 9030 13897 9058 13902
rect 8526 13790 8834 13818
rect 8526 13593 8554 13790
rect 8526 13567 8527 13593
rect 8553 13567 8554 13593
rect 8526 13561 8554 13567
rect 7462 13435 7490 13454
rect 8414 13426 8498 13454
rect 8134 12866 8162 12871
rect 8134 12819 8162 12838
rect 8022 12810 8050 12815
rect 7126 12385 7154 12390
rect 7910 12641 7938 12647
rect 7910 12615 7911 12641
rect 7937 12615 7938 12641
rect 7910 12418 7938 12615
rect 7910 12385 7938 12390
rect 6398 12361 6482 12362
rect 6398 12335 6455 12361
rect 6481 12335 6482 12361
rect 6398 12334 6482 12335
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 4998 12026 5026 12031
rect 4998 11979 5026 11998
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 6398 11970 6426 12334
rect 6454 12329 6482 12334
rect 7966 12362 7994 12367
rect 6846 12306 6874 12311
rect 6846 12259 6874 12278
rect 7910 12306 7938 12311
rect 7966 12306 7994 12334
rect 7910 12305 7994 12306
rect 7910 12279 7911 12305
rect 7937 12279 7994 12305
rect 7910 12278 7994 12279
rect 7910 12273 7938 12278
rect 6958 12026 6986 12031
rect 6398 11923 6426 11942
rect 6734 11970 6762 11975
rect 6062 11914 6090 11919
rect 6062 11913 6258 11914
rect 6062 11887 6063 11913
rect 6089 11887 6258 11913
rect 6062 11886 6258 11887
rect 6062 11881 6090 11886
rect 6230 11689 6258 11886
rect 6230 11663 6231 11689
rect 6257 11663 6258 11689
rect 6230 11657 6258 11663
rect 6734 11858 6762 11942
rect 6790 11858 6818 11863
rect 6734 11857 6818 11858
rect 6734 11831 6791 11857
rect 6817 11831 6818 11857
rect 6734 11830 6818 11831
rect 6286 11578 6314 11583
rect 6286 11531 6314 11550
rect 2086 11489 2114 11494
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 6342 11130 6370 11135
rect 6342 11083 6370 11102
rect 6174 11074 6202 11079
rect 5894 11073 6202 11074
rect 5894 11047 6175 11073
rect 6201 11047 6202 11073
rect 5894 11046 6202 11047
rect 5894 10849 5922 11046
rect 6174 11041 6202 11046
rect 5894 10823 5895 10849
rect 5921 10823 5922 10849
rect 5894 10817 5922 10823
rect 5558 10794 5586 10799
rect 6734 10794 6762 11830
rect 6790 11825 6818 11830
rect 6846 11690 6874 11695
rect 6846 11633 6874 11662
rect 6846 11607 6847 11633
rect 6873 11607 6874 11633
rect 6846 11601 6874 11607
rect 6902 11633 6930 11639
rect 6902 11607 6903 11633
rect 6929 11607 6930 11633
rect 6790 11130 6818 11135
rect 6790 11083 6818 11102
rect 6790 10794 6818 10799
rect 6734 10766 6790 10794
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 5558 10094 5586 10766
rect 6790 10761 6818 10766
rect 6902 10094 6930 11607
rect 6958 11633 6986 11998
rect 7854 12026 7882 12031
rect 7854 11969 7882 11998
rect 7854 11943 7855 11969
rect 7881 11943 7882 11969
rect 7854 11937 7882 11943
rect 7686 11857 7714 11863
rect 7686 11831 7687 11857
rect 7713 11831 7714 11857
rect 7182 11690 7210 11695
rect 7126 11662 7182 11690
rect 6958 11607 6959 11633
rect 6985 11607 6986 11633
rect 6958 11601 6986 11607
rect 7070 11634 7098 11639
rect 7070 11587 7098 11606
rect 7014 11578 7042 11583
rect 7014 11531 7042 11550
rect 7070 11242 7098 11247
rect 7126 11242 7154 11662
rect 7182 11643 7210 11662
rect 7294 11689 7322 11695
rect 7294 11663 7295 11689
rect 7321 11663 7322 11689
rect 7238 11634 7266 11639
rect 7294 11634 7322 11663
rect 7266 11606 7322 11634
rect 7238 11601 7266 11606
rect 7070 11241 7154 11242
rect 7070 11215 7071 11241
rect 7097 11215 7154 11241
rect 7070 11214 7154 11215
rect 7070 11209 7098 11214
rect 6958 11186 6986 11191
rect 6958 11139 6986 11158
rect 7294 11018 7322 11606
rect 7350 11634 7378 11639
rect 7350 11587 7378 11606
rect 7686 11634 7714 11831
rect 7798 11858 7826 11863
rect 7798 11811 7826 11830
rect 8022 11857 8050 12782
rect 8190 12754 8218 12759
rect 8022 11831 8023 11857
rect 8049 11831 8050 11857
rect 7686 11601 7714 11606
rect 7294 10985 7322 10990
rect 7854 10962 7882 10967
rect 7854 10849 7882 10934
rect 7854 10823 7855 10849
rect 7881 10823 7882 10849
rect 7854 10817 7882 10823
rect 7182 10794 7210 10799
rect 7182 10747 7210 10766
rect 7462 10794 7490 10799
rect 6958 10737 6986 10743
rect 6958 10711 6959 10737
rect 6985 10711 6986 10737
rect 6958 10458 6986 10711
rect 7294 10458 7322 10463
rect 6958 10457 7322 10458
rect 6958 10431 7295 10457
rect 7321 10431 7322 10457
rect 6958 10430 7322 10431
rect 6958 10401 6986 10430
rect 7294 10425 7322 10430
rect 7462 10458 7490 10766
rect 7574 10794 7602 10799
rect 8022 10794 8050 11831
rect 8078 12726 8190 12754
rect 8078 11970 8106 12726
rect 8190 12707 8218 12726
rect 8078 10905 8106 11942
rect 8134 12641 8162 12647
rect 8134 12615 8135 12641
rect 8161 12615 8162 12641
rect 8134 11634 8162 12615
rect 8302 12642 8330 12647
rect 8246 12417 8274 12423
rect 8246 12391 8247 12417
rect 8273 12391 8274 12417
rect 8246 12306 8274 12391
rect 8302 12362 8330 12614
rect 8358 12641 8386 12647
rect 8358 12615 8359 12641
rect 8385 12615 8386 12641
rect 8358 12474 8386 12615
rect 8358 12441 8386 12446
rect 8358 12362 8386 12367
rect 8302 12361 8386 12362
rect 8302 12335 8359 12361
rect 8385 12335 8386 12361
rect 8302 12334 8386 12335
rect 8358 12329 8386 12334
rect 8190 12026 8218 12031
rect 8190 11979 8218 11998
rect 8246 11914 8274 12278
rect 8414 12026 8442 13426
rect 8638 13202 8666 13790
rect 8806 13594 8834 13599
rect 8694 13538 8722 13543
rect 8694 13481 8722 13510
rect 8806 13537 8834 13566
rect 9198 13593 9226 13902
rect 9422 13874 9450 13879
rect 10486 13874 10514 15946
rect 12110 14377 12138 15946
rect 12110 14351 12111 14377
rect 12137 14351 12138 14377
rect 10710 14322 10738 14327
rect 11046 14322 11074 14327
rect 10710 14275 10738 14294
rect 10878 14321 11074 14322
rect 10878 14295 11047 14321
rect 11073 14295 11074 14321
rect 10878 14294 11074 14295
rect 10878 14041 10906 14294
rect 11046 14289 11074 14294
rect 10878 14015 10879 14041
rect 10905 14015 10906 14041
rect 10878 14009 10906 14015
rect 11438 14266 11466 14271
rect 9422 13873 9562 13874
rect 9422 13847 9423 13873
rect 9449 13847 9562 13873
rect 9422 13846 9562 13847
rect 9422 13841 9450 13846
rect 9198 13567 9199 13593
rect 9225 13567 9226 13593
rect 9198 13561 9226 13567
rect 9534 13593 9562 13846
rect 10374 13873 10514 13874
rect 10374 13847 10487 13873
rect 10513 13847 10514 13873
rect 10374 13846 10514 13847
rect 9534 13567 9535 13593
rect 9561 13567 9562 13593
rect 9534 13561 9562 13567
rect 9590 13594 9618 13599
rect 8806 13511 8807 13537
rect 8833 13511 8834 13537
rect 8806 13505 8834 13511
rect 8918 13537 8946 13543
rect 8918 13511 8919 13537
rect 8945 13511 8946 13537
rect 8694 13455 8695 13481
rect 8721 13455 8722 13481
rect 8694 13314 8722 13455
rect 8750 13482 8778 13487
rect 8918 13454 8946 13511
rect 9478 13538 9506 13543
rect 9478 13491 9506 13510
rect 9590 13537 9618 13566
rect 9590 13511 9591 13537
rect 9617 13511 9618 13537
rect 9590 13505 9618 13511
rect 9814 13538 9842 13543
rect 10094 13538 10122 13543
rect 9814 13537 10122 13538
rect 9814 13511 9815 13537
rect 9841 13511 10095 13537
rect 10121 13511 10122 13537
rect 9814 13510 10122 13511
rect 9814 13505 9842 13510
rect 10094 13505 10122 13510
rect 10374 13537 10402 13846
rect 10486 13841 10514 13846
rect 10710 13985 10738 13991
rect 10710 13959 10711 13985
rect 10737 13959 10738 13985
rect 10374 13511 10375 13537
rect 10401 13511 10402 13537
rect 10374 13505 10402 13511
rect 8750 13435 8778 13454
rect 8862 13426 8946 13454
rect 10150 13482 10178 13487
rect 10150 13481 10234 13482
rect 10150 13455 10151 13481
rect 10177 13455 10234 13481
rect 10150 13454 10234 13455
rect 10150 13449 10178 13454
rect 9702 13426 9730 13431
rect 10038 13426 10066 13431
rect 10206 13426 10290 13454
rect 8694 13286 8778 13314
rect 8694 13202 8722 13207
rect 8638 13201 8722 13202
rect 8638 13175 8695 13201
rect 8721 13175 8722 13201
rect 8638 13174 8722 13175
rect 8694 13169 8722 13174
rect 8750 13146 8778 13286
rect 8862 13257 8890 13426
rect 9702 13425 9842 13426
rect 9702 13399 9703 13425
rect 9729 13399 9842 13425
rect 9702 13398 9842 13399
rect 9702 13393 9730 13398
rect 8862 13231 8863 13257
rect 8889 13231 8890 13257
rect 8862 13225 8890 13231
rect 8806 13146 8834 13151
rect 8750 13145 8834 13146
rect 8750 13119 8807 13145
rect 8833 13119 8834 13145
rect 8750 13118 8834 13119
rect 8806 12866 8834 13118
rect 8806 12833 8834 12838
rect 8918 13145 8946 13151
rect 8918 13119 8919 13145
rect 8945 13119 8946 13145
rect 8918 12698 8946 13119
rect 8974 13145 9002 13151
rect 8974 13119 8975 13145
rect 9001 13119 9002 13145
rect 8974 12754 9002 13119
rect 9814 13034 9842 13398
rect 10038 13425 10122 13426
rect 10038 13399 10039 13425
rect 10065 13399 10122 13425
rect 10038 13398 10122 13399
rect 10038 13393 10066 13398
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10094 13258 10122 13398
rect 10038 13230 10122 13258
rect 9814 13006 9954 13034
rect 9926 12865 9954 13006
rect 9926 12839 9927 12865
rect 9953 12839 9954 12865
rect 9926 12833 9954 12839
rect 9030 12810 9058 12815
rect 9030 12763 9058 12782
rect 8974 12721 9002 12726
rect 9870 12698 9898 12703
rect 8862 12670 8918 12698
rect 8526 12641 8554 12647
rect 8526 12615 8527 12641
rect 8553 12615 8554 12641
rect 8526 12362 8554 12615
rect 8526 12329 8554 12334
rect 8750 12474 8778 12479
rect 8750 12250 8778 12446
rect 8862 12473 8890 12670
rect 8918 12651 8946 12670
rect 9590 12697 9898 12698
rect 9590 12671 9871 12697
rect 9897 12671 9898 12697
rect 9590 12670 9898 12671
rect 8974 12642 9002 12647
rect 8974 12595 9002 12614
rect 8862 12447 8863 12473
rect 8889 12447 8890 12473
rect 8862 12441 8890 12447
rect 8918 12417 8946 12423
rect 8918 12391 8919 12417
rect 8945 12391 8946 12417
rect 8806 12250 8834 12255
rect 8750 12249 8834 12250
rect 8750 12223 8807 12249
rect 8833 12223 8834 12249
rect 8750 12222 8834 12223
rect 8750 12026 8778 12222
rect 8806 12217 8834 12222
rect 8414 12025 8498 12026
rect 8414 11999 8415 12025
rect 8441 11999 8498 12025
rect 8414 11998 8498 11999
rect 8414 11993 8442 11998
rect 8246 11881 8274 11886
rect 8302 11969 8330 11975
rect 8302 11943 8303 11969
rect 8329 11943 8330 11969
rect 8302 11802 8330 11943
rect 8302 11769 8330 11774
rect 8134 11601 8162 11606
rect 8414 11633 8442 11639
rect 8414 11607 8415 11633
rect 8441 11607 8442 11633
rect 8302 11578 8330 11583
rect 8078 10879 8079 10905
rect 8105 10879 8106 10905
rect 8078 10873 8106 10879
rect 8134 11185 8162 11191
rect 8134 11159 8135 11185
rect 8161 11159 8162 11185
rect 8134 10794 8162 11159
rect 8302 10962 8330 11550
rect 8414 11466 8442 11607
rect 8358 11438 8414 11466
rect 8358 11185 8386 11438
rect 8414 11433 8442 11438
rect 8358 11159 8359 11185
rect 8385 11159 8386 11185
rect 8358 11153 8386 11159
rect 8414 11186 8442 11191
rect 8470 11186 8498 11998
rect 8526 11970 8554 11975
rect 8526 11923 8554 11942
rect 8582 11913 8610 11919
rect 8582 11887 8583 11913
rect 8609 11887 8610 11913
rect 8582 11858 8610 11887
rect 8582 11690 8610 11830
rect 8582 11657 8610 11662
rect 8638 11802 8666 11807
rect 8470 11158 8554 11186
rect 8414 11139 8442 11158
rect 7574 10793 7658 10794
rect 7574 10767 7575 10793
rect 7601 10767 7658 10793
rect 7574 10766 7658 10767
rect 8022 10766 8162 10794
rect 7574 10761 7602 10766
rect 6958 10375 6959 10401
rect 6985 10375 6986 10401
rect 6958 10369 6986 10375
rect 7406 10401 7434 10407
rect 7406 10375 7407 10401
rect 7433 10375 7434 10401
rect 7126 10289 7154 10295
rect 7126 10263 7127 10289
rect 7153 10263 7154 10289
rect 7126 10234 7154 10263
rect 7126 10201 7154 10206
rect 5558 10066 5754 10094
rect 6902 10066 7098 10094
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 5726 9225 5754 10066
rect 7070 10065 7154 10066
rect 7070 10039 7071 10065
rect 7097 10039 7154 10065
rect 7070 10038 7154 10039
rect 7070 10033 7098 10038
rect 5726 9199 5727 9225
rect 5753 9199 5754 9225
rect 5726 9193 5754 9199
rect 6118 9506 6146 9511
rect 6118 9225 6146 9478
rect 6118 9199 6119 9225
rect 6145 9199 6146 9225
rect 6118 9193 6146 9199
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5726 8834 5754 8839
rect 7126 8834 7154 10038
rect 7238 10009 7266 10015
rect 7238 9983 7239 10009
rect 7265 9983 7266 10009
rect 7238 9954 7266 9983
rect 7238 9921 7266 9926
rect 7406 10010 7434 10375
rect 7406 9786 7434 9982
rect 7182 9758 7434 9786
rect 7182 9169 7210 9758
rect 7182 9143 7183 9169
rect 7209 9143 7210 9169
rect 7182 9137 7210 9143
rect 7406 9226 7434 9231
rect 7462 9226 7490 10430
rect 7574 10290 7602 10295
rect 7574 10243 7602 10262
rect 7630 10234 7658 10766
rect 7854 10458 7882 10463
rect 7854 10411 7882 10430
rect 7630 10201 7658 10206
rect 7910 10010 7938 10015
rect 7910 9963 7938 9982
rect 7630 9954 7658 9959
rect 7630 9907 7658 9926
rect 8134 9730 8162 10766
rect 8246 10794 8274 10799
rect 8302 10794 8330 10934
rect 8470 11073 8498 11079
rect 8470 11047 8471 11073
rect 8497 11047 8498 11073
rect 8470 10850 8498 11047
rect 8470 10817 8498 10822
rect 8246 10793 8330 10794
rect 8246 10767 8247 10793
rect 8273 10767 8330 10793
rect 8246 10766 8330 10767
rect 8358 10793 8386 10799
rect 8358 10767 8359 10793
rect 8385 10767 8386 10793
rect 8246 10761 8274 10766
rect 8358 10122 8386 10767
rect 8190 10094 8386 10122
rect 8190 10009 8218 10094
rect 8190 9983 8191 10009
rect 8217 9983 8218 10009
rect 8190 9977 8218 9983
rect 8246 10010 8274 10015
rect 8190 9730 8218 9735
rect 8134 9702 8190 9730
rect 8190 9697 8218 9702
rect 8246 9617 8274 9982
rect 8358 10010 8386 10094
rect 8358 9977 8386 9982
rect 8358 9674 8386 9679
rect 8358 9627 8386 9646
rect 8246 9591 8247 9617
rect 8273 9591 8274 9617
rect 8246 9585 8274 9591
rect 8526 9618 8554 11158
rect 8638 10066 8666 11774
rect 8694 11634 8722 11639
rect 8694 10793 8722 11606
rect 8750 10962 8778 11998
rect 8918 11970 8946 12391
rect 8918 11802 8946 11942
rect 8974 12306 9002 12311
rect 8974 11913 9002 12278
rect 9422 12306 9450 12311
rect 9422 12259 9450 12278
rect 9590 12026 9618 12670
rect 9870 12665 9898 12670
rect 9926 12642 9954 12661
rect 10038 12642 10066 13230
rect 10038 12614 10122 12642
rect 9926 12609 9954 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10094 12474 10122 12614
rect 10038 12446 10122 12474
rect 9646 12362 9674 12367
rect 9646 12315 9674 12334
rect 9422 12025 9618 12026
rect 9422 11999 9591 12025
rect 9617 11999 9618 12025
rect 9422 11998 9618 11999
rect 9366 11970 9394 11975
rect 8974 11887 8975 11913
rect 9001 11887 9002 11913
rect 8974 11881 9002 11887
rect 9198 11969 9394 11970
rect 9198 11943 9367 11969
rect 9393 11943 9394 11969
rect 9198 11942 9394 11943
rect 8918 11769 8946 11774
rect 9030 11633 9058 11639
rect 9030 11607 9031 11633
rect 9057 11607 9058 11633
rect 8862 11578 8890 11583
rect 8974 11578 9002 11583
rect 8890 11577 9002 11578
rect 8890 11551 8975 11577
rect 9001 11551 9002 11577
rect 8890 11550 9002 11551
rect 8806 11522 8834 11527
rect 8806 11475 8834 11494
rect 8806 11186 8834 11191
rect 8862 11186 8890 11550
rect 8974 11545 9002 11550
rect 8806 11185 8890 11186
rect 8806 11159 8807 11185
rect 8833 11159 8890 11185
rect 8806 11158 8890 11159
rect 8806 11153 8834 11158
rect 9030 11130 9058 11607
rect 8974 11129 9058 11130
rect 8974 11103 9031 11129
rect 9057 11103 9058 11129
rect 8974 11102 9058 11103
rect 8750 10934 8890 10962
rect 8694 10767 8695 10793
rect 8721 10767 8722 10793
rect 8694 10761 8722 10767
rect 8694 10066 8722 10071
rect 8638 10065 8722 10066
rect 8638 10039 8695 10065
rect 8721 10039 8722 10065
rect 8638 10038 8722 10039
rect 8694 10033 8722 10038
rect 8862 9953 8890 10934
rect 8862 9927 8863 9953
rect 8889 9927 8890 9953
rect 8862 9921 8890 9927
rect 8918 10850 8946 10855
rect 8806 9730 8834 9735
rect 8638 9618 8666 9623
rect 8526 9617 8610 9618
rect 8526 9591 8527 9617
rect 8553 9591 8610 9617
rect 8526 9590 8610 9591
rect 8526 9585 8554 9590
rect 7406 9225 7490 9226
rect 7406 9199 7407 9225
rect 7433 9199 7490 9225
rect 7406 9198 7490 9199
rect 8470 9338 8498 9343
rect 7294 8834 7322 8839
rect 7126 8833 7322 8834
rect 7126 8807 7295 8833
rect 7321 8807 7322 8833
rect 7126 8806 7322 8807
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 5726 8385 5754 8806
rect 6790 8666 6818 8671
rect 6790 8497 6818 8638
rect 6790 8471 6791 8497
rect 6817 8471 6818 8497
rect 6790 8465 6818 8471
rect 7182 8610 7210 8615
rect 5726 8359 5727 8385
rect 5753 8359 5754 8385
rect 5726 8353 5754 8359
rect 5838 8442 5866 8447
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8073 994 8078
rect 1022 8105 1050 8111
rect 1022 8079 1023 8105
rect 1049 8079 1050 8105
rect 1022 7770 1050 8079
rect 2142 8050 2170 8055
rect 2142 8003 2170 8022
rect 1022 7737 1050 7742
rect 5838 7601 5866 8414
rect 7182 8441 7210 8582
rect 7182 8415 7183 8441
rect 7209 8415 7210 8441
rect 6902 8386 6930 8391
rect 5838 7575 5839 7601
rect 5865 7575 5866 7601
rect 5838 7569 5866 7575
rect 5894 8050 5922 8055
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 5894 6817 5922 8022
rect 6902 7713 6930 8358
rect 6902 7687 6903 7713
rect 6929 7687 6930 7713
rect 6902 7681 6930 7687
rect 6958 7938 6986 7943
rect 6958 6929 6986 7910
rect 7182 7658 7210 8415
rect 7294 8498 7322 8806
rect 7350 8834 7378 8839
rect 7350 8777 7378 8806
rect 7350 8751 7351 8777
rect 7377 8751 7378 8777
rect 7350 8745 7378 8751
rect 7406 8610 7434 9198
rect 7966 8890 7994 8895
rect 7686 8833 7714 8839
rect 7686 8807 7687 8833
rect 7713 8807 7714 8833
rect 7462 8722 7490 8727
rect 7462 8675 7490 8694
rect 7406 8577 7434 8582
rect 7350 8498 7378 8503
rect 7294 8497 7378 8498
rect 7294 8471 7351 8497
rect 7377 8471 7378 8497
rect 7294 8470 7378 8471
rect 7238 8050 7266 8055
rect 7294 8050 7322 8470
rect 7350 8465 7378 8470
rect 7406 8498 7434 8503
rect 7406 8451 7434 8470
rect 7518 8442 7546 8447
rect 7518 8395 7546 8414
rect 7686 8442 7714 8807
rect 7854 8834 7882 8839
rect 7854 8787 7882 8806
rect 7966 8833 7994 8862
rect 7966 8807 7967 8833
rect 7993 8807 7994 8833
rect 7742 8722 7770 8727
rect 7742 8675 7770 8694
rect 7798 8721 7826 8727
rect 7798 8695 7799 8721
rect 7825 8695 7826 8721
rect 7798 8666 7826 8695
rect 7798 8633 7826 8638
rect 7966 8553 7994 8807
rect 8470 8889 8498 9310
rect 8582 8945 8610 9590
rect 8638 9226 8666 9590
rect 8806 9617 8834 9702
rect 8806 9591 8807 9617
rect 8833 9591 8834 9617
rect 8806 9585 8834 9591
rect 8918 9618 8946 10822
rect 8918 9585 8946 9590
rect 8974 9674 9002 11102
rect 9030 11097 9058 11102
rect 9142 11298 9170 11303
rect 9142 11018 9170 11270
rect 9142 10794 9170 10990
rect 9086 10793 9170 10794
rect 9086 10767 9143 10793
rect 9169 10767 9170 10793
rect 9086 10766 9170 10767
rect 9086 9898 9114 10766
rect 9142 10761 9170 10766
rect 9198 10905 9226 11942
rect 9366 11937 9394 11942
rect 9198 10879 9199 10905
rect 9225 10879 9226 10905
rect 9086 9865 9114 9870
rect 9142 10290 9170 10295
rect 8694 9505 8722 9511
rect 8694 9479 8695 9505
rect 8721 9479 8722 9505
rect 8694 9338 8722 9479
rect 8750 9506 8778 9511
rect 8750 9459 8778 9478
rect 8694 9310 8778 9338
rect 8694 9226 8722 9231
rect 8638 9225 8722 9226
rect 8638 9199 8695 9225
rect 8721 9199 8722 9225
rect 8638 9198 8722 9199
rect 8694 9193 8722 9198
rect 8582 8919 8583 8945
rect 8609 8919 8610 8945
rect 8582 8913 8610 8919
rect 8470 8863 8471 8889
rect 8497 8863 8498 8889
rect 8470 8834 8498 8863
rect 8750 8834 8778 9310
rect 8974 9225 9002 9646
rect 9142 9674 9170 10262
rect 9142 9627 9170 9646
rect 8974 9199 8975 9225
rect 9001 9199 9002 9225
rect 8974 9193 9002 9199
rect 9086 9618 9114 9623
rect 8918 8834 8946 8839
rect 8750 8806 8918 8834
rect 8470 8801 8498 8806
rect 8918 8777 8946 8806
rect 9086 8833 9114 9590
rect 9086 8807 9087 8833
rect 9113 8807 9114 8833
rect 9086 8801 9114 8807
rect 8918 8751 8919 8777
rect 8945 8751 8946 8777
rect 8918 8745 8946 8751
rect 8750 8722 8778 8727
rect 8750 8721 8890 8722
rect 8750 8695 8751 8721
rect 8777 8695 8890 8721
rect 8750 8694 8890 8695
rect 8750 8689 8778 8694
rect 7966 8527 7967 8553
rect 7993 8527 7994 8553
rect 7966 8521 7994 8527
rect 8246 8610 8274 8615
rect 8246 8553 8274 8582
rect 8246 8527 8247 8553
rect 8273 8527 8274 8553
rect 8246 8521 8274 8527
rect 7742 8442 7770 8447
rect 7686 8441 7770 8442
rect 7686 8415 7743 8441
rect 7769 8415 7770 8441
rect 7686 8414 7770 8415
rect 7238 8049 7322 8050
rect 7238 8023 7239 8049
rect 7265 8023 7322 8049
rect 7238 8022 7322 8023
rect 7350 8050 7378 8055
rect 7238 8017 7266 8022
rect 7294 7938 7322 7943
rect 7350 7938 7378 8022
rect 7686 8049 7714 8414
rect 7742 8330 7770 8414
rect 7798 8442 7826 8447
rect 7798 8395 7826 8414
rect 7910 8442 7938 8447
rect 7910 8395 7938 8414
rect 7854 8386 7882 8391
rect 7854 8339 7882 8358
rect 7742 8297 7770 8302
rect 7686 8023 7687 8049
rect 7713 8023 7714 8049
rect 7686 8017 7714 8023
rect 7798 8106 7826 8111
rect 7798 8049 7826 8078
rect 8862 8106 8890 8694
rect 9142 8442 9170 8447
rect 9198 8442 9226 10879
rect 9254 10066 9282 10071
rect 9254 9617 9282 10038
rect 9366 10010 9394 10015
rect 9366 9963 9394 9982
rect 9254 9591 9255 9617
rect 9281 9591 9282 9617
rect 9254 9585 9282 9591
rect 9310 9898 9338 9903
rect 9254 9338 9282 9343
rect 9310 9338 9338 9870
rect 9422 9674 9450 11998
rect 9590 11993 9618 11998
rect 9982 11969 10010 11975
rect 9982 11943 9983 11969
rect 10009 11943 10010 11969
rect 9814 11914 9842 11919
rect 9814 11867 9842 11886
rect 9758 11857 9786 11863
rect 9758 11831 9759 11857
rect 9785 11831 9786 11857
rect 9590 11522 9618 11527
rect 9590 10793 9618 11494
rect 9590 10767 9591 10793
rect 9617 10767 9618 10793
rect 9590 10761 9618 10767
rect 9646 11185 9674 11191
rect 9646 11159 9647 11185
rect 9673 11159 9674 11185
rect 9478 10234 9506 10239
rect 9478 10010 9506 10206
rect 9646 10066 9674 11159
rect 9646 10033 9674 10038
rect 9478 10009 9618 10010
rect 9478 9983 9479 10009
rect 9505 9983 9618 10009
rect 9478 9982 9618 9983
rect 9478 9977 9506 9982
rect 9254 9337 9338 9338
rect 9254 9311 9255 9337
rect 9281 9311 9338 9337
rect 9254 9310 9338 9311
rect 9366 9673 9450 9674
rect 9366 9647 9423 9673
rect 9449 9647 9450 9673
rect 9366 9646 9450 9647
rect 9254 9305 9282 9310
rect 9254 8890 9282 8895
rect 9254 8843 9282 8862
rect 9310 8778 9338 8783
rect 9366 8778 9394 9646
rect 9422 9641 9450 9646
rect 9534 9897 9562 9903
rect 9534 9871 9535 9897
rect 9561 9871 9562 9897
rect 9422 9562 9450 9567
rect 9422 9226 9450 9534
rect 9534 9338 9562 9871
rect 9590 9562 9618 9982
rect 9702 9954 9730 9959
rect 9702 9618 9730 9926
rect 9758 9730 9786 11831
rect 9982 11858 10010 11943
rect 10038 11858 10066 12446
rect 10262 12418 10290 13426
rect 10710 12865 10738 13959
rect 11270 13986 11298 13991
rect 11270 13939 11298 13958
rect 10822 13930 10850 13935
rect 10934 13930 10962 13935
rect 10822 13883 10850 13902
rect 10878 13929 10962 13930
rect 10878 13903 10935 13929
rect 10961 13903 10962 13929
rect 10878 13902 10962 13903
rect 10878 13594 10906 13902
rect 10934 13897 10962 13902
rect 11214 13930 11242 13935
rect 11214 13883 11242 13902
rect 10878 13257 10906 13566
rect 11438 13537 11466 14238
rect 12110 13986 12138 14351
rect 12334 14322 12362 14327
rect 12334 14275 12362 14294
rect 12110 13953 12138 13958
rect 12894 13594 12922 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 20118 17345 20146 17351
rect 20118 17319 20119 17345
rect 20145 17319 20146 17345
rect 20118 17178 20146 17319
rect 20118 17145 20146 17150
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 11438 13511 11439 13537
rect 11465 13511 11466 13537
rect 11046 13314 11074 13319
rect 10878 13231 10879 13257
rect 10905 13231 10906 13257
rect 10878 13225 10906 13231
rect 10990 13286 11046 13314
rect 10710 12839 10711 12865
rect 10737 12839 10738 12865
rect 10710 12833 10738 12839
rect 10990 12753 11018 13286
rect 11046 13281 11074 13286
rect 11438 13314 11466 13511
rect 12670 13593 12922 13594
rect 12670 13567 12895 13593
rect 12921 13567 12922 13593
rect 12670 13566 12922 13567
rect 11830 13482 11858 13487
rect 11438 13281 11466 13286
rect 11606 13481 11858 13482
rect 11606 13455 11831 13481
rect 11857 13455 11858 13481
rect 11606 13454 11858 13455
rect 11606 13257 11634 13454
rect 11830 13449 11858 13454
rect 11606 13231 11607 13257
rect 11633 13231 11634 13257
rect 11606 13225 11634 13231
rect 11158 13174 11522 13202
rect 11046 13146 11074 13151
rect 11158 13146 11186 13174
rect 11046 13145 11186 13146
rect 11046 13119 11047 13145
rect 11073 13119 11186 13145
rect 11046 13118 11186 13119
rect 11494 13146 11522 13174
rect 12670 13201 12698 13566
rect 12894 13561 12922 13566
rect 13118 13425 13146 13431
rect 13118 13399 13119 13425
rect 13145 13399 13146 13425
rect 12670 13175 12671 13201
rect 12697 13175 12698 13201
rect 12670 13169 12698 13175
rect 12726 13314 12754 13319
rect 11550 13146 11578 13151
rect 11494 13145 11578 13146
rect 11494 13119 11551 13145
rect 11577 13119 11578 13145
rect 11494 13118 11578 13119
rect 11046 13113 11074 13118
rect 11438 13089 11466 13095
rect 11438 13063 11439 13089
rect 11465 13063 11466 13089
rect 11214 13034 11242 13039
rect 11214 13033 11298 13034
rect 11214 13007 11215 13033
rect 11241 13007 11298 13033
rect 11214 13006 11298 13007
rect 11214 13001 11242 13006
rect 10990 12727 10991 12753
rect 11017 12727 11018 12753
rect 10990 12721 11018 12727
rect 10654 12698 10682 12703
rect 10654 12651 10682 12670
rect 10262 12371 10290 12390
rect 10710 12641 10738 12647
rect 10710 12615 10711 12641
rect 10737 12615 10738 12641
rect 10150 12362 10178 12367
rect 10150 12026 10178 12334
rect 10710 12194 10738 12615
rect 10710 12161 10738 12166
rect 10822 12306 10850 12311
rect 10150 11993 10178 11998
rect 10654 12026 10682 12031
rect 10654 11979 10682 11998
rect 9982 11830 10122 11858
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9814 11689 9842 11695
rect 9814 11663 9815 11689
rect 9841 11663 9842 11689
rect 9814 9842 9842 11663
rect 10094 11186 10122 11830
rect 10206 11857 10234 11863
rect 10206 11831 10207 11857
rect 10233 11831 10234 11857
rect 10206 11298 10234 11831
rect 10374 11858 10402 11863
rect 10374 11811 10402 11830
rect 10710 11858 10738 11863
rect 10710 11857 10794 11858
rect 10710 11831 10711 11857
rect 10737 11831 10794 11857
rect 10710 11830 10794 11831
rect 10710 11825 10738 11830
rect 10262 11690 10290 11695
rect 10262 11633 10290 11662
rect 10262 11607 10263 11633
rect 10289 11607 10290 11633
rect 10262 11601 10290 11607
rect 10206 11270 10290 11298
rect 10262 11242 10290 11270
rect 10206 11186 10234 11191
rect 10094 11158 10206 11186
rect 10206 11129 10234 11158
rect 10206 11103 10207 11129
rect 10233 11103 10234 11129
rect 10206 11097 10234 11103
rect 9926 11074 9954 11093
rect 9926 11041 9954 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10206 10962 10234 10967
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10206 10121 10234 10934
rect 10206 10095 10207 10121
rect 10233 10095 10234 10121
rect 10206 10089 10234 10095
rect 9982 10066 10010 10071
rect 9982 9953 10010 10038
rect 10262 10010 10290 11214
rect 10710 11130 10738 11135
rect 10710 11083 10738 11102
rect 10262 9977 10290 9982
rect 10374 11073 10402 11079
rect 10374 11047 10375 11073
rect 10401 11047 10402 11073
rect 9982 9927 9983 9953
rect 10009 9927 10010 9953
rect 9982 9921 10010 9927
rect 9814 9814 10066 9842
rect 9870 9730 9898 9735
rect 9758 9702 9842 9730
rect 9758 9618 9786 9623
rect 9702 9617 9786 9618
rect 9702 9591 9759 9617
rect 9785 9591 9786 9617
rect 9702 9590 9786 9591
rect 9758 9585 9786 9590
rect 9590 9534 9730 9562
rect 9534 9305 9562 9310
rect 9646 9450 9674 9455
rect 9422 9225 9618 9226
rect 9422 9199 9423 9225
rect 9449 9199 9618 9225
rect 9422 9198 9618 9199
rect 9422 9193 9450 9198
rect 9422 9114 9450 9119
rect 9422 8945 9450 9086
rect 9422 8919 9423 8945
rect 9449 8919 9450 8945
rect 9422 8913 9450 8919
rect 9590 8889 9618 9198
rect 9590 8863 9591 8889
rect 9617 8863 9618 8889
rect 9590 8857 9618 8863
rect 9310 8777 9394 8778
rect 9310 8751 9311 8777
rect 9337 8751 9394 8777
rect 9310 8750 9394 8751
rect 9310 8745 9338 8750
rect 9142 8441 9226 8442
rect 9142 8415 9143 8441
rect 9169 8415 9226 8441
rect 9142 8414 9226 8415
rect 9254 8497 9282 8503
rect 9254 8471 9255 8497
rect 9281 8471 9282 8497
rect 8890 8078 9002 8106
rect 8862 8059 8890 8078
rect 7798 8023 7799 8049
rect 7825 8023 7826 8049
rect 7798 8017 7826 8023
rect 7406 7994 7434 7999
rect 7518 7994 7546 7999
rect 7406 7993 7546 7994
rect 7406 7967 7407 7993
rect 7433 7967 7519 7993
rect 7545 7967 7546 7993
rect 7406 7966 7546 7967
rect 7406 7961 7434 7966
rect 7518 7961 7546 7966
rect 7294 7937 7378 7938
rect 7294 7911 7295 7937
rect 7321 7911 7378 7937
rect 7294 7910 7378 7911
rect 7574 7938 7602 7943
rect 8918 7938 8946 7943
rect 7294 7905 7322 7910
rect 7574 7891 7602 7910
rect 8750 7937 8946 7938
rect 8750 7911 8919 7937
rect 8945 7911 8946 7937
rect 8750 7910 8946 7911
rect 7238 7658 7266 7663
rect 7518 7658 7546 7663
rect 7182 7657 7546 7658
rect 7182 7631 7239 7657
rect 7265 7631 7519 7657
rect 7545 7631 7546 7657
rect 7182 7630 7546 7631
rect 7238 7625 7266 7630
rect 7406 7266 7434 7630
rect 7518 7625 7546 7630
rect 7742 7602 7770 7607
rect 7742 7321 7770 7574
rect 7742 7295 7743 7321
rect 7769 7295 7770 7321
rect 7742 7289 7770 7295
rect 6958 6903 6959 6929
rect 6985 6903 6986 6929
rect 6958 6897 6986 6903
rect 7350 7265 7602 7266
rect 7350 7239 7407 7265
rect 7433 7239 7602 7265
rect 7350 7238 7602 7239
rect 7350 6873 7378 7238
rect 7406 7233 7434 7238
rect 7574 7154 7602 7238
rect 7574 6985 7602 7126
rect 7574 6959 7575 6985
rect 7601 6959 7602 6985
rect 7574 6953 7602 6959
rect 8750 7154 8778 7910
rect 8918 7905 8946 7910
rect 8806 7714 8834 7719
rect 8806 7667 8834 7686
rect 8918 7658 8946 7663
rect 8974 7658 9002 8078
rect 9142 7770 9170 8414
rect 9254 8386 9282 8471
rect 9254 8353 9282 8358
rect 9142 7742 9338 7770
rect 9142 7713 9170 7742
rect 9142 7687 9143 7713
rect 9169 7687 9170 7713
rect 9142 7681 9170 7687
rect 9254 7658 9282 7663
rect 8918 7657 9002 7658
rect 8918 7631 8919 7657
rect 8945 7631 9002 7657
rect 8918 7630 9002 7631
rect 9198 7657 9282 7658
rect 9198 7631 9255 7657
rect 9281 7631 9282 7657
rect 9198 7630 9282 7631
rect 8918 7625 8946 7630
rect 8862 7602 8890 7621
rect 9198 7574 9226 7630
rect 9254 7625 9282 7630
rect 8862 7569 8890 7574
rect 9030 7545 9058 7551
rect 9030 7519 9031 7545
rect 9057 7519 9058 7545
rect 9030 7490 9058 7519
rect 9030 7457 9058 7462
rect 9086 7546 9226 7574
rect 9030 7378 9058 7383
rect 9086 7378 9114 7546
rect 9198 7490 9226 7495
rect 9198 7434 9226 7462
rect 9198 7406 9282 7434
rect 9030 7377 9114 7378
rect 9030 7351 9031 7377
rect 9057 7351 9114 7377
rect 9030 7350 9114 7351
rect 9030 7345 9058 7350
rect 8806 7321 8834 7327
rect 9198 7322 9226 7327
rect 8806 7295 8807 7321
rect 8833 7295 8834 7321
rect 8806 7210 8834 7295
rect 9086 7321 9226 7322
rect 9086 7295 9199 7321
rect 9225 7295 9226 7321
rect 9086 7294 9226 7295
rect 8974 7210 9002 7215
rect 8806 7209 9002 7210
rect 8806 7183 8975 7209
rect 9001 7183 9002 7209
rect 8806 7182 9002 7183
rect 7350 6847 7351 6873
rect 7377 6847 7378 6873
rect 7350 6841 7378 6847
rect 8750 6874 8778 7126
rect 8750 6873 8834 6874
rect 8750 6847 8751 6873
rect 8777 6847 8834 6873
rect 8750 6846 8834 6847
rect 8750 6841 8778 6846
rect 5894 6791 5895 6817
rect 5921 6791 5922 6817
rect 5894 6785 5922 6791
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 8806 6538 8834 6846
rect 8806 6537 8946 6538
rect 8806 6511 8807 6537
rect 8833 6511 8946 6537
rect 8806 6510 8946 6511
rect 8806 6505 8834 6510
rect 8918 6481 8946 6510
rect 8918 6455 8919 6481
rect 8945 6455 8946 6481
rect 8918 6449 8946 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8974 2169 9002 7182
rect 9086 6929 9114 7294
rect 9198 7289 9226 7294
rect 9254 7210 9282 7406
rect 9310 7210 9338 7742
rect 9646 7378 9674 9422
rect 9702 8834 9730 9534
rect 9814 8946 9842 9702
rect 9870 9673 9898 9702
rect 9870 9647 9871 9673
rect 9897 9647 9898 9673
rect 9870 9641 9898 9647
rect 9870 9561 9898 9567
rect 9870 9535 9871 9561
rect 9897 9535 9898 9561
rect 9870 9506 9898 9535
rect 10038 9506 10066 9814
rect 10374 9674 10402 11047
rect 10654 11074 10682 11079
rect 10654 10514 10682 11046
rect 10710 10962 10738 10967
rect 10766 10962 10794 11830
rect 10738 10934 10794 10962
rect 10822 11577 10850 12278
rect 11102 12194 11130 12199
rect 11130 12166 11186 12194
rect 11102 12161 11130 12166
rect 11046 11970 11074 11989
rect 11046 11937 11074 11942
rect 10822 11551 10823 11577
rect 10849 11551 10850 11577
rect 10822 10962 10850 11551
rect 11046 11857 11074 11863
rect 11046 11831 11047 11857
rect 11073 11831 11074 11857
rect 10878 11074 10906 11079
rect 10878 11027 10906 11046
rect 11046 11074 11074 11831
rect 11158 11690 11186 12166
rect 11158 11643 11186 11662
rect 11214 11858 11242 11863
rect 11102 11633 11130 11639
rect 11102 11607 11103 11633
rect 11129 11607 11130 11633
rect 11102 11298 11130 11607
rect 11214 11633 11242 11830
rect 11214 11607 11215 11633
rect 11241 11607 11242 11633
rect 11214 11601 11242 11607
rect 11102 11265 11130 11270
rect 11158 11186 11186 11191
rect 11046 11041 11074 11046
rect 11102 11185 11186 11186
rect 11102 11159 11159 11185
rect 11185 11159 11186 11185
rect 11102 11158 11186 11159
rect 10822 10934 10906 10962
rect 10710 10929 10738 10934
rect 10822 10738 10850 10743
rect 10654 10486 10794 10514
rect 10654 10401 10682 10407
rect 10654 10375 10655 10401
rect 10681 10375 10682 10401
rect 10654 10234 10682 10375
rect 10430 10206 10682 10234
rect 10430 10065 10458 10206
rect 10430 10039 10431 10065
rect 10457 10039 10458 10065
rect 10430 9954 10458 10039
rect 10430 9921 10458 9926
rect 10486 10121 10514 10127
rect 10486 10095 10487 10121
rect 10513 10095 10514 10121
rect 10374 9641 10402 9646
rect 10318 9617 10346 9623
rect 10318 9591 10319 9617
rect 10345 9591 10346 9617
rect 10318 9506 10346 9591
rect 10038 9478 10178 9506
rect 9870 9473 9898 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10150 9226 10178 9478
rect 10150 9193 10178 9198
rect 10206 9478 10318 9506
rect 9814 8918 10010 8946
rect 9702 8833 9786 8834
rect 9702 8807 9703 8833
rect 9729 8807 9786 8833
rect 9702 8806 9786 8807
rect 9702 8801 9730 8806
rect 9758 8778 9786 8806
rect 9926 8833 9954 8839
rect 9926 8807 9927 8833
rect 9953 8807 9954 8833
rect 9926 8778 9954 8807
rect 9758 8750 9954 8778
rect 9982 8722 10010 8918
rect 10206 8889 10234 9478
rect 10318 9473 10346 9478
rect 10486 9282 10514 10095
rect 10710 9618 10738 9623
rect 10710 9571 10738 9590
rect 10486 9235 10514 9254
rect 10654 9338 10682 9343
rect 10206 8863 10207 8889
rect 10233 8863 10234 8889
rect 10206 8857 10234 8863
rect 10654 8889 10682 9310
rect 10766 9225 10794 10486
rect 10822 10289 10850 10710
rect 10822 10263 10823 10289
rect 10849 10263 10850 10289
rect 10822 10257 10850 10263
rect 10878 10345 10906 10934
rect 10878 10319 10879 10345
rect 10905 10319 10906 10345
rect 10878 10122 10906 10319
rect 10878 10089 10906 10094
rect 10990 10345 11018 10351
rect 10990 10319 10991 10345
rect 11017 10319 11018 10345
rect 10934 9730 10962 9735
rect 10934 9617 10962 9702
rect 10934 9591 10935 9617
rect 10961 9591 10962 9617
rect 10934 9585 10962 9591
rect 10990 9506 11018 10319
rect 11102 10010 11130 11158
rect 11158 11153 11186 11158
rect 11214 11186 11242 11191
rect 11270 11186 11298 13006
rect 11326 13033 11354 13039
rect 11326 13007 11327 13033
rect 11353 13007 11354 13033
rect 11326 12418 11354 13007
rect 11382 12698 11410 12703
rect 11438 12698 11466 13063
rect 11382 12697 11466 12698
rect 11382 12671 11383 12697
rect 11409 12671 11466 12697
rect 11382 12670 11466 12671
rect 11382 12665 11410 12670
rect 11326 11354 11354 12390
rect 11438 12642 11466 12670
rect 11382 12305 11410 12311
rect 11382 12279 11383 12305
rect 11409 12279 11410 12305
rect 11382 11970 11410 12279
rect 11382 11937 11410 11942
rect 11382 11802 11410 11807
rect 11382 11466 11410 11774
rect 11438 11746 11466 12614
rect 11438 11713 11466 11718
rect 11494 11858 11522 11863
rect 11438 11633 11466 11639
rect 11438 11607 11439 11633
rect 11465 11607 11466 11633
rect 11438 11578 11466 11607
rect 11438 11545 11466 11550
rect 11494 11633 11522 11830
rect 11550 11802 11578 13118
rect 11662 13146 11690 13151
rect 11662 13099 11690 13118
rect 12614 13146 12642 13151
rect 12614 13099 12642 13118
rect 12446 12809 12474 12815
rect 12446 12783 12447 12809
rect 12473 12783 12474 12809
rect 11662 12474 11690 12479
rect 11662 12427 11690 12446
rect 12110 12474 12138 12479
rect 12110 12427 12138 12446
rect 12446 12474 12474 12783
rect 12670 12810 12698 12815
rect 12726 12810 12754 13286
rect 13118 13314 13146 13399
rect 13118 13281 13146 13286
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 12670 12809 12866 12810
rect 12670 12783 12671 12809
rect 12697 12783 12866 12809
rect 12670 12782 12866 12783
rect 12670 12777 12698 12782
rect 12446 12441 12474 12446
rect 11550 11769 11578 11774
rect 11886 12305 11914 12311
rect 11886 12279 11887 12305
rect 11913 12279 11914 12305
rect 11494 11607 11495 11633
rect 11521 11607 11522 11633
rect 11438 11466 11466 11471
rect 11382 11465 11466 11466
rect 11382 11439 11439 11465
rect 11465 11439 11466 11465
rect 11382 11438 11466 11439
rect 11494 11466 11522 11607
rect 11662 11746 11690 11751
rect 11494 11438 11634 11466
rect 11438 11433 11466 11438
rect 11326 11326 11466 11354
rect 11382 11242 11410 11247
rect 11382 11195 11410 11214
rect 11242 11158 11298 11186
rect 11326 11185 11354 11191
rect 11326 11159 11327 11185
rect 11353 11159 11354 11185
rect 11214 11153 11242 11158
rect 11214 11073 11242 11079
rect 11214 11047 11215 11073
rect 11241 11047 11242 11073
rect 11158 10737 11186 10743
rect 11158 10711 11159 10737
rect 11185 10711 11186 10737
rect 11158 10402 11186 10711
rect 11158 10355 11186 10374
rect 11158 10010 11186 10015
rect 11102 10009 11186 10010
rect 11102 9983 11159 10009
rect 11185 9983 11186 10009
rect 11102 9982 11186 9983
rect 11102 9562 11130 9982
rect 11158 9977 11186 9982
rect 11102 9529 11130 9534
rect 11158 9617 11186 9623
rect 11158 9591 11159 9617
rect 11185 9591 11186 9617
rect 10990 9473 11018 9478
rect 11158 9506 11186 9591
rect 11158 9473 11186 9478
rect 11102 9282 11130 9287
rect 10766 9199 10767 9225
rect 10793 9199 10794 9225
rect 10766 8946 10794 9199
rect 10934 9226 10962 9231
rect 10934 9179 10962 9198
rect 10766 8913 10794 8918
rect 10654 8863 10655 8889
rect 10681 8863 10682 8889
rect 10654 8857 10682 8863
rect 10710 8834 10738 8839
rect 10822 8834 10850 8839
rect 10710 8833 10822 8834
rect 10710 8807 10711 8833
rect 10737 8807 10822 8833
rect 10710 8806 10822 8807
rect 10710 8801 10738 8806
rect 10822 8787 10850 8806
rect 11102 8833 11130 9254
rect 11102 8807 11103 8833
rect 11129 8807 11130 8833
rect 11102 8801 11130 8807
rect 11046 8777 11074 8783
rect 11046 8751 11047 8777
rect 11073 8751 11074 8777
rect 9646 7345 9674 7350
rect 9814 8694 10010 8722
rect 10934 8721 10962 8727
rect 10934 8695 10935 8721
rect 10961 8695 10962 8721
rect 9366 7322 9394 7327
rect 9590 7322 9618 7327
rect 9366 7321 9618 7322
rect 9366 7295 9367 7321
rect 9393 7295 9591 7321
rect 9617 7295 9618 7321
rect 9366 7294 9618 7295
rect 9366 7289 9394 7294
rect 9590 7289 9618 7294
rect 9814 7322 9842 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10654 8554 10682 8559
rect 10934 8554 10962 8695
rect 10654 8507 10682 8526
rect 10766 8526 10962 8554
rect 10710 8385 10738 8391
rect 10710 8359 10711 8385
rect 10737 8359 10738 8385
rect 10710 7938 10738 8359
rect 10766 8385 10794 8526
rect 10766 8359 10767 8385
rect 10793 8359 10794 8385
rect 10766 8353 10794 8359
rect 10878 8442 10906 8447
rect 10710 7905 10738 7910
rect 10822 7994 10850 7999
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9926 7602 9954 7621
rect 9926 7569 9954 7574
rect 10822 7602 10850 7966
rect 9982 7378 10010 7383
rect 9982 7331 10010 7350
rect 9814 7289 9842 7294
rect 10150 7322 10178 7327
rect 10430 7322 10458 7327
rect 10150 7321 10346 7322
rect 10150 7295 10151 7321
rect 10177 7295 10346 7321
rect 10150 7294 10346 7295
rect 10150 7289 10178 7294
rect 9758 7266 9786 7271
rect 9758 7219 9786 7238
rect 9534 7210 9562 7215
rect 9310 7209 9562 7210
rect 9310 7183 9535 7209
rect 9561 7183 9562 7209
rect 9310 7182 9562 7183
rect 9254 7163 9282 7182
rect 9534 7177 9562 7182
rect 9702 7209 9730 7215
rect 9702 7183 9703 7209
rect 9729 7183 9730 7209
rect 9086 6903 9087 6929
rect 9113 6903 9114 6929
rect 9086 6897 9114 6903
rect 9702 6818 9730 7183
rect 10094 7153 10122 7159
rect 10094 7127 10095 7153
rect 10121 7127 10122 7153
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9814 6818 9842 6823
rect 9702 6790 9814 6818
rect 9310 6762 9338 6767
rect 9310 6537 9338 6734
rect 9310 6511 9311 6537
rect 9337 6511 9338 6537
rect 9310 6505 9338 6511
rect 8974 2143 8975 2169
rect 9001 2143 9002 2169
rect 8974 2137 9002 2143
rect 8750 2058 8778 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8750 400 8778 2030
rect 9254 2058 9282 2063
rect 9254 2011 9282 2030
rect 9814 1778 9842 6790
rect 10094 6538 10122 7127
rect 10318 6873 10346 7294
rect 10374 7154 10402 7159
rect 10374 7107 10402 7126
rect 10318 6847 10319 6873
rect 10345 6847 10346 6873
rect 10318 6841 10346 6847
rect 10430 6873 10458 7294
rect 10430 6847 10431 6873
rect 10457 6847 10458 6873
rect 10430 6841 10458 6847
rect 10542 7210 10570 7215
rect 10542 6873 10570 7182
rect 10542 6847 10543 6873
rect 10569 6847 10570 6873
rect 10542 6841 10570 6847
rect 10150 6818 10178 6823
rect 10150 6771 10178 6790
rect 10598 6762 10626 6767
rect 10598 6715 10626 6734
rect 10374 6538 10402 6543
rect 10094 6537 10402 6538
rect 10094 6511 10375 6537
rect 10401 6511 10402 6537
rect 10094 6510 10402 6511
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10374 2169 10402 6510
rect 10374 2143 10375 2169
rect 10401 2143 10402 2169
rect 10374 2137 10402 2143
rect 10094 2058 10122 2063
rect 9870 1778 9898 1783
rect 9814 1777 9898 1778
rect 9814 1751 9871 1777
rect 9897 1751 9898 1777
rect 9814 1750 9898 1751
rect 9870 1745 9898 1750
rect 9590 1666 9618 1671
rect 9590 1665 9786 1666
rect 9590 1639 9591 1665
rect 9617 1639 9786 1665
rect 9590 1638 9786 1639
rect 9590 1633 9618 1638
rect 9758 400 9786 1638
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10094 400 10122 2030
rect 10710 2058 10738 2063
rect 10710 2011 10738 2030
rect 10822 1777 10850 7574
rect 10878 7377 10906 8414
rect 11046 7994 11074 8751
rect 11214 8554 11242 11047
rect 11326 10962 11354 11159
rect 11326 10929 11354 10934
rect 11382 10122 11410 10127
rect 11382 10009 11410 10094
rect 11382 9983 11383 10009
rect 11409 9983 11410 10009
rect 11382 9977 11410 9983
rect 11438 9730 11466 11326
rect 11606 10682 11634 11438
rect 11662 11130 11690 11718
rect 11830 11690 11858 11695
rect 11718 11633 11746 11639
rect 11718 11607 11719 11633
rect 11745 11607 11746 11633
rect 11718 11242 11746 11607
rect 11718 11209 11746 11214
rect 11830 11241 11858 11662
rect 11886 11634 11914 12279
rect 11886 11587 11914 11606
rect 12110 11914 12138 11919
rect 12110 11577 12138 11886
rect 12390 11858 12418 11863
rect 12110 11551 12111 11577
rect 12137 11551 12138 11577
rect 12110 11297 12138 11551
rect 12110 11271 12111 11297
rect 12137 11271 12138 11297
rect 12110 11265 12138 11271
rect 12222 11577 12250 11583
rect 12222 11551 12223 11577
rect 12249 11551 12250 11577
rect 11830 11215 11831 11241
rect 11857 11215 11858 11241
rect 11830 11209 11858 11215
rect 11662 11097 11690 11102
rect 11942 11185 11970 11191
rect 11942 11159 11943 11185
rect 11969 11159 11970 11185
rect 11942 11018 11970 11159
rect 11942 10985 11970 10990
rect 12166 11074 12194 11079
rect 11606 10649 11634 10654
rect 12110 10066 12138 10071
rect 12166 10066 12194 11046
rect 12222 10178 12250 11551
rect 12390 11577 12418 11830
rect 12390 11551 12391 11577
rect 12417 11551 12418 11577
rect 12390 11545 12418 11551
rect 12838 11577 12866 12782
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 13062 12026 13090 12031
rect 13062 12025 13202 12026
rect 13062 11999 13063 12025
rect 13089 11999 13202 12025
rect 13062 11998 13202 11999
rect 13062 11993 13090 11998
rect 12894 11914 12922 11919
rect 12894 11867 12922 11886
rect 13006 11858 13034 11863
rect 12838 11551 12839 11577
rect 12865 11551 12866 11577
rect 12278 11522 12306 11527
rect 12278 11475 12306 11494
rect 12838 11354 12866 11551
rect 12838 11321 12866 11326
rect 12950 11857 13034 11858
rect 12950 11831 13007 11857
rect 13033 11831 13034 11857
rect 12950 11830 13034 11831
rect 12502 11242 12530 11247
rect 12950 11242 12978 11830
rect 13006 11825 13034 11830
rect 12278 11186 12306 11191
rect 12278 11139 12306 11158
rect 12390 11186 12418 11191
rect 12390 11185 12474 11186
rect 12390 11159 12391 11185
rect 12417 11159 12474 11185
rect 12390 11158 12474 11159
rect 12390 11153 12418 11158
rect 12334 11074 12362 11079
rect 12334 11073 12418 11074
rect 12334 11047 12335 11073
rect 12361 11047 12418 11073
rect 12334 11046 12418 11047
rect 12334 11041 12362 11046
rect 12222 10150 12362 10178
rect 12278 10066 12306 10071
rect 12166 10065 12306 10066
rect 12166 10039 12279 10065
rect 12305 10039 12306 10065
rect 12166 10038 12306 10039
rect 11438 9697 11466 9702
rect 11494 9729 11522 9735
rect 11494 9703 11495 9729
rect 11521 9703 11522 9729
rect 11326 9618 11354 9623
rect 11326 9571 11354 9590
rect 11382 9617 11410 9623
rect 11382 9591 11383 9617
rect 11409 9591 11410 9617
rect 11046 7961 11074 7966
rect 11102 8526 11214 8554
rect 10990 7938 11018 7943
rect 10990 7713 11018 7910
rect 10990 7687 10991 7713
rect 11017 7687 11018 7713
rect 10990 7681 11018 7687
rect 10878 7351 10879 7377
rect 10905 7351 10906 7377
rect 10878 7345 10906 7351
rect 11046 7322 11074 7327
rect 11046 7275 11074 7294
rect 11102 7266 11130 8526
rect 11214 8521 11242 8526
rect 11270 9337 11298 9343
rect 11270 9311 11271 9337
rect 11297 9311 11298 9337
rect 11270 7490 11298 9311
rect 11382 9338 11410 9591
rect 11382 9305 11410 9310
rect 11438 9282 11466 9287
rect 11438 8889 11466 9254
rect 11494 9281 11522 9703
rect 11718 9674 11746 9679
rect 11718 9627 11746 9646
rect 12110 9673 12138 10038
rect 12110 9647 12111 9673
rect 12137 9647 12138 9673
rect 12110 9641 12138 9647
rect 11494 9255 11495 9281
rect 11521 9255 11522 9281
rect 11494 9249 11522 9255
rect 11662 9562 11690 9567
rect 11494 8946 11522 8951
rect 11494 8899 11522 8918
rect 11438 8863 11439 8889
rect 11465 8863 11466 8889
rect 11438 8857 11466 8863
rect 11326 8834 11354 8839
rect 11326 8787 11354 8806
rect 11550 8554 11578 8559
rect 11550 8161 11578 8526
rect 11550 8135 11551 8161
rect 11577 8135 11578 8161
rect 11550 8129 11578 8135
rect 11662 8105 11690 9534
rect 12278 9561 12306 10038
rect 12278 9535 12279 9561
rect 12305 9535 12306 9561
rect 12278 9529 12306 9535
rect 12334 9506 12362 10150
rect 12390 10122 12418 11046
rect 12390 10089 12418 10094
rect 12446 10066 12474 11158
rect 12502 11185 12530 11214
rect 12502 11159 12503 11185
rect 12529 11159 12530 11185
rect 12502 11130 12530 11159
rect 12782 11214 12978 11242
rect 13006 11354 13034 11359
rect 12502 11102 12698 11130
rect 12614 10793 12642 10799
rect 12614 10767 12615 10793
rect 12641 10767 12642 10793
rect 12614 10346 12642 10767
rect 12558 10318 12642 10346
rect 12670 10794 12698 11102
rect 12782 10905 12810 11214
rect 13006 11186 13034 11326
rect 13174 11242 13202 11998
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 13286 11970 13314 11975
rect 13230 11913 13258 11919
rect 13230 11887 13231 11913
rect 13257 11887 13258 11913
rect 13230 11634 13258 11887
rect 13286 11913 13314 11942
rect 13958 11970 13986 11975
rect 13958 11923 13986 11942
rect 14294 11970 14322 11975
rect 13286 11887 13287 11913
rect 13313 11887 13314 11913
rect 13286 11881 13314 11887
rect 13398 11858 13426 11863
rect 13398 11811 13426 11830
rect 14070 11858 14098 11863
rect 14070 11811 14098 11830
rect 13230 11606 13314 11634
rect 13230 11522 13258 11527
rect 13230 11475 13258 11494
rect 13230 11242 13258 11247
rect 13174 11241 13258 11242
rect 13174 11215 13231 11241
rect 13257 11215 13258 11241
rect 13174 11214 13258 11215
rect 13230 11209 13258 11214
rect 12894 11179 13034 11186
rect 12894 11153 12895 11179
rect 12921 11158 13034 11179
rect 12921 11153 12922 11158
rect 12894 11147 12922 11153
rect 13006 11018 13034 11158
rect 12782 10879 12783 10905
rect 12809 10879 12810 10905
rect 12782 10873 12810 10879
rect 12838 10906 12866 10911
rect 12838 10859 12866 10878
rect 12950 10850 12978 10855
rect 12950 10803 12978 10822
rect 12726 10794 12754 10799
rect 12670 10793 12754 10794
rect 12670 10767 12727 10793
rect 12753 10767 12754 10793
rect 12670 10766 12754 10767
rect 12558 10066 12586 10318
rect 12446 10033 12474 10038
rect 12502 10038 12586 10066
rect 12446 9618 12474 9623
rect 12502 9618 12530 10038
rect 12474 9590 12530 9618
rect 12614 9618 12642 9623
rect 12670 9618 12698 10766
rect 12726 10761 12754 10766
rect 12950 10682 12978 10687
rect 12614 9617 12698 9618
rect 12614 9591 12615 9617
rect 12641 9591 12698 9617
rect 12614 9590 12698 9591
rect 12726 10122 12754 10127
rect 12726 9617 12754 10094
rect 12950 9618 12978 10654
rect 13006 10457 13034 10990
rect 13062 11130 13090 11135
rect 13286 11130 13314 11606
rect 13062 10626 13090 11102
rect 13174 11102 13314 11130
rect 13902 11578 13930 11583
rect 13174 10906 13202 11102
rect 13174 10859 13202 10878
rect 13398 11018 13426 11023
rect 13118 10738 13146 10743
rect 13118 10691 13146 10710
rect 13062 10598 13146 10626
rect 13006 10431 13007 10457
rect 13033 10431 13034 10457
rect 13006 10425 13034 10431
rect 12726 9591 12727 9617
rect 12753 9591 12754 9617
rect 12446 9571 12474 9590
rect 12614 9562 12642 9590
rect 12726 9585 12754 9591
rect 12782 9617 12978 9618
rect 12782 9591 12951 9617
rect 12977 9591 12978 9617
rect 12782 9590 12978 9591
rect 12614 9529 12642 9534
rect 12558 9506 12586 9511
rect 12782 9506 12810 9590
rect 12950 9585 12978 9590
rect 13062 9730 13090 9735
rect 13062 9617 13090 9702
rect 13062 9591 13063 9617
rect 13089 9591 13090 9617
rect 13062 9585 13090 9591
rect 13006 9506 13034 9511
rect 12334 9505 12586 9506
rect 12334 9479 12559 9505
rect 12585 9479 12586 9505
rect 12334 9478 12586 9479
rect 12166 9282 12194 9287
rect 12166 9235 12194 9254
rect 12278 9282 12306 9287
rect 12334 9282 12362 9478
rect 12558 9473 12586 9478
rect 12726 9478 12810 9506
rect 12894 9505 13034 9506
rect 12894 9479 13007 9505
rect 13033 9479 13034 9505
rect 12894 9478 13034 9479
rect 12278 9281 12362 9282
rect 12278 9255 12279 9281
rect 12305 9255 12362 9281
rect 12278 9254 12362 9255
rect 12670 9281 12698 9287
rect 12670 9255 12671 9281
rect 12697 9255 12698 9281
rect 12278 9249 12306 9254
rect 11718 9226 11746 9231
rect 11718 8833 11746 9198
rect 11998 9225 12026 9231
rect 11998 9199 11999 9225
rect 12025 9199 12026 9225
rect 11998 9170 12026 9199
rect 11998 9137 12026 9142
rect 12054 9225 12082 9231
rect 12054 9199 12055 9225
rect 12081 9199 12082 9225
rect 12054 9002 12082 9199
rect 12558 9225 12586 9231
rect 12558 9199 12559 9225
rect 12585 9199 12586 9225
rect 11718 8807 11719 8833
rect 11745 8807 11746 8833
rect 11718 8801 11746 8807
rect 11998 8974 12082 9002
rect 12110 9169 12138 9175
rect 12110 9143 12111 9169
rect 12137 9143 12138 9169
rect 11998 8386 12026 8974
rect 12054 8890 12082 8895
rect 12110 8890 12138 9143
rect 12558 9170 12586 9199
rect 12558 9137 12586 9142
rect 12670 9114 12698 9255
rect 12726 9281 12754 9478
rect 12894 9338 12922 9478
rect 13006 9473 13034 9478
rect 13118 9394 13146 10598
rect 13174 9506 13202 9511
rect 13174 9459 13202 9478
rect 13398 9506 13426 10990
rect 13902 10094 13930 11550
rect 14294 11521 14322 11942
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 18830 11858 18858 11863
rect 18830 11577 18858 11830
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 18830 11551 18831 11577
rect 18857 11551 18858 11577
rect 18830 11545 18858 11551
rect 14294 11495 14295 11521
rect 14321 11495 14322 11521
rect 14294 11489 14322 11495
rect 14518 11521 14546 11527
rect 14518 11495 14519 11521
rect 14545 11495 14546 11521
rect 14294 11242 14322 11247
rect 14294 10850 14322 11214
rect 14518 11242 14546 11495
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 14630 11242 14658 11247
rect 14518 11241 14658 11242
rect 14518 11215 14631 11241
rect 14657 11215 14658 11241
rect 14518 11214 14658 11215
rect 14518 11018 14546 11214
rect 14630 11209 14658 11214
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 14518 10985 14546 10990
rect 14294 10817 14322 10822
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 13790 10066 13930 10094
rect 18942 10401 18970 10407
rect 18942 10375 18943 10401
rect 18969 10375 18970 10401
rect 13622 9561 13650 9567
rect 13622 9535 13623 9561
rect 13649 9535 13650 9561
rect 13454 9506 13482 9511
rect 13398 9505 13482 9506
rect 13398 9479 13455 9505
rect 13481 9479 13482 9505
rect 13398 9478 13482 9479
rect 12726 9255 12727 9281
rect 12753 9255 12754 9281
rect 12726 9249 12754 9255
rect 12782 9310 12922 9338
rect 13006 9366 13146 9394
rect 13006 9337 13034 9366
rect 13006 9311 13007 9337
rect 13033 9311 13034 9337
rect 12670 9081 12698 9086
rect 12054 8889 12138 8890
rect 12054 8863 12055 8889
rect 12081 8863 12138 8889
rect 12054 8862 12138 8863
rect 12054 8857 12082 8862
rect 12782 8442 12810 9310
rect 13006 9305 13034 9311
rect 12950 9282 12978 9287
rect 12894 9281 12978 9282
rect 12894 9255 12951 9281
rect 12977 9255 12978 9281
rect 12894 9254 12978 9255
rect 12782 8409 12810 8414
rect 12838 9226 12866 9231
rect 12838 8554 12866 9198
rect 12894 8946 12922 9254
rect 12950 9249 12978 9254
rect 13118 9226 13146 9231
rect 13398 9226 13426 9478
rect 13454 9473 13482 9478
rect 13118 9225 13202 9226
rect 13118 9199 13119 9225
rect 13145 9199 13202 9225
rect 13118 9198 13202 9199
rect 13118 9193 13146 9198
rect 12894 8913 12922 8918
rect 13118 9114 13146 9119
rect 13118 8889 13146 9086
rect 13118 8863 13119 8889
rect 13145 8863 13146 8889
rect 13118 8857 13146 8863
rect 13174 8834 13202 9198
rect 13230 8834 13258 8839
rect 13174 8833 13258 8834
rect 13174 8807 13231 8833
rect 13257 8807 13258 8833
rect 13174 8806 13258 8807
rect 12838 8553 13034 8554
rect 12838 8527 12839 8553
rect 12865 8527 13034 8553
rect 12838 8526 13034 8527
rect 11998 8353 12026 8358
rect 11662 8079 11663 8105
rect 11689 8079 11690 8105
rect 11662 8073 11690 8079
rect 11382 7938 11410 7943
rect 11382 7937 11746 7938
rect 11382 7911 11383 7937
rect 11409 7911 11746 7937
rect 11382 7910 11746 7911
rect 11382 7905 11410 7910
rect 11382 7657 11410 7663
rect 11382 7631 11383 7657
rect 11409 7631 11410 7657
rect 11382 7602 11410 7631
rect 11606 7602 11634 7607
rect 11382 7601 11634 7602
rect 11382 7575 11607 7601
rect 11633 7575 11634 7601
rect 11382 7546 11634 7575
rect 11718 7574 11746 7910
rect 12838 7657 12866 8526
rect 13006 8441 13034 8526
rect 13006 8415 13007 8441
rect 13033 8415 13034 8441
rect 13006 8409 13034 8415
rect 13230 7714 13258 8806
rect 13342 8721 13370 8727
rect 13342 8695 13343 8721
rect 13369 8695 13370 8721
rect 13342 8498 13370 8695
rect 13398 8722 13426 9198
rect 13622 9114 13650 9535
rect 13734 9562 13762 9567
rect 13734 9515 13762 9534
rect 13790 9450 13818 10066
rect 18830 10010 18858 10015
rect 18774 10009 18858 10010
rect 18774 9983 18831 10009
rect 18857 9983 18858 10009
rect 18774 9982 18858 9983
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 13846 9674 13874 9679
rect 14070 9674 14098 9679
rect 13846 9673 14098 9674
rect 13846 9647 13847 9673
rect 13873 9647 14071 9673
rect 14097 9647 14098 9673
rect 13846 9646 14098 9647
rect 13846 9641 13874 9646
rect 14070 9641 14098 9646
rect 14686 9617 14714 9623
rect 14686 9591 14687 9617
rect 14713 9591 14714 9617
rect 13902 9561 13930 9567
rect 13902 9535 13903 9561
rect 13929 9535 13930 9561
rect 13902 9450 13930 9535
rect 14686 9562 14714 9591
rect 14686 9529 14714 9534
rect 14798 9618 14826 9623
rect 14798 9561 14826 9590
rect 15022 9617 15050 9623
rect 15022 9591 15023 9617
rect 15049 9591 15050 9617
rect 14798 9535 14799 9561
rect 14825 9535 14826 9561
rect 14798 9529 14826 9535
rect 14854 9562 14882 9567
rect 14126 9506 14154 9511
rect 13622 9081 13650 9086
rect 13734 9422 13930 9450
rect 13958 9505 14154 9506
rect 13958 9479 14127 9505
rect 14153 9479 14154 9505
rect 13958 9478 14154 9479
rect 13510 8890 13538 8895
rect 13510 8833 13538 8862
rect 13510 8807 13511 8833
rect 13537 8807 13538 8833
rect 13454 8778 13482 8783
rect 13454 8731 13482 8750
rect 13398 8689 13426 8694
rect 13398 8498 13426 8503
rect 13342 8497 13426 8498
rect 13342 8471 13399 8497
rect 13425 8471 13426 8497
rect 13342 8470 13426 8471
rect 13398 8465 13426 8470
rect 13510 8162 13538 8807
rect 13734 8833 13762 9422
rect 13958 9338 13986 9478
rect 14126 9473 14154 9478
rect 14182 9505 14210 9511
rect 14182 9479 14183 9505
rect 14209 9479 14210 9505
rect 13790 9310 13986 9338
rect 13790 9281 13818 9310
rect 13790 9255 13791 9281
rect 13817 9255 13818 9281
rect 13790 9249 13818 9255
rect 14182 8890 14210 9479
rect 14854 9169 14882 9534
rect 15022 9562 15050 9591
rect 15022 9529 15050 9534
rect 15134 9506 15162 9511
rect 15134 9459 15162 9478
rect 18774 9506 18802 9982
rect 18830 9977 18858 9982
rect 18942 9730 18970 10375
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 18942 9697 18970 9702
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 18774 9473 18802 9478
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 18830 9226 18858 9231
rect 18830 9179 18858 9198
rect 14854 9143 14855 9169
rect 14881 9143 14882 9169
rect 14854 9137 14882 9143
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 14182 8857 14210 8862
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 13734 8807 13735 8833
rect 13761 8807 13762 8833
rect 13734 8801 13762 8807
rect 13790 8834 13818 8839
rect 13790 8777 13818 8806
rect 14462 8834 14490 8839
rect 13790 8751 13791 8777
rect 13817 8751 13818 8777
rect 13790 8745 13818 8751
rect 13902 8778 13930 8783
rect 13902 8731 13930 8750
rect 14070 8722 14098 8727
rect 14070 8675 14098 8694
rect 14462 8385 14490 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 14462 8359 14463 8385
rect 14489 8359 14490 8385
rect 14462 8353 14490 8359
rect 14518 8722 14546 8727
rect 13566 8162 13594 8167
rect 13510 8161 13594 8162
rect 13510 8135 13567 8161
rect 13593 8135 13594 8161
rect 13510 8134 13594 8135
rect 13566 8129 13594 8134
rect 13734 8050 13762 8055
rect 13734 8003 13762 8022
rect 14294 8050 14322 8055
rect 13230 7681 13258 7686
rect 13622 7937 13650 7943
rect 13622 7911 13623 7937
rect 13649 7911 13650 7937
rect 12838 7631 12839 7657
rect 12865 7631 12866 7657
rect 11718 7546 11802 7574
rect 11270 7462 11466 7490
rect 11438 7434 11466 7462
rect 11438 7377 11466 7406
rect 11438 7351 11439 7377
rect 11465 7351 11466 7377
rect 11438 7345 11466 7351
rect 11382 7322 11410 7327
rect 11382 7275 11410 7294
rect 11102 7233 11130 7238
rect 11270 7266 11298 7271
rect 11270 7219 11298 7238
rect 11214 7209 11242 7215
rect 11214 7183 11215 7209
rect 11241 7183 11242 7209
rect 10990 7153 11018 7159
rect 10990 7127 10991 7153
rect 11017 7127 11018 7153
rect 10878 6874 10906 6879
rect 10878 6827 10906 6846
rect 10990 6818 11018 7127
rect 11214 6929 11242 7183
rect 11214 6903 11215 6929
rect 11241 6903 11242 6929
rect 11214 6897 11242 6903
rect 11438 7154 11466 7159
rect 11438 6874 11466 7126
rect 11606 7154 11634 7546
rect 11718 7434 11746 7439
rect 11718 7377 11746 7406
rect 11718 7351 11719 7377
rect 11745 7351 11746 7377
rect 11718 7345 11746 7351
rect 11774 7266 11802 7546
rect 12614 7378 12642 7383
rect 11830 7266 11858 7271
rect 11774 7265 11858 7266
rect 11774 7239 11831 7265
rect 11857 7239 11858 7265
rect 11774 7238 11858 7239
rect 11606 7121 11634 7126
rect 11662 7209 11690 7215
rect 11662 7183 11663 7209
rect 11689 7183 11690 7209
rect 11046 6818 11074 6823
rect 10990 6790 11046 6818
rect 11046 6785 11074 6790
rect 11438 6481 11466 6846
rect 11662 6538 11690 7183
rect 11718 7210 11746 7215
rect 11774 7210 11802 7238
rect 11830 7233 11858 7238
rect 11942 7266 11970 7271
rect 11942 7219 11970 7238
rect 11746 7182 11802 7210
rect 11718 7177 11746 7182
rect 12390 7154 12418 7159
rect 12390 7107 12418 7126
rect 12614 6929 12642 7350
rect 12670 7266 12698 7271
rect 12670 6985 12698 7238
rect 12838 7154 12866 7631
rect 13230 7601 13258 7607
rect 13622 7602 13650 7911
rect 13230 7575 13231 7601
rect 13257 7575 13258 7601
rect 13174 7378 13202 7383
rect 13174 7265 13202 7350
rect 13230 7321 13258 7575
rect 13342 7574 13650 7602
rect 14294 7601 14322 8022
rect 14518 7769 14546 8694
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 18830 8050 18858 8055
rect 18830 8003 18858 8022
rect 14518 7743 14519 7769
rect 14545 7743 14546 7769
rect 14518 7737 14546 7743
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 14294 7575 14295 7601
rect 14321 7575 14322 7601
rect 13342 7377 13370 7574
rect 14294 7569 14322 7575
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13342 7351 13343 7377
rect 13369 7351 13370 7377
rect 13342 7345 13370 7351
rect 13230 7295 13231 7321
rect 13257 7295 13258 7321
rect 13230 7289 13258 7295
rect 13174 7239 13175 7265
rect 13201 7239 13202 7265
rect 13174 7233 13202 7239
rect 12838 7121 12866 7126
rect 13118 7154 13146 7159
rect 12670 6959 12671 6985
rect 12697 6959 12698 6985
rect 12670 6953 12698 6959
rect 12614 6903 12615 6929
rect 12641 6903 12642 6929
rect 12614 6897 12642 6903
rect 12782 6874 12810 6879
rect 12782 6873 12866 6874
rect 12782 6847 12783 6873
rect 12809 6847 12866 6873
rect 12782 6846 12866 6847
rect 12782 6841 12810 6846
rect 12278 6818 12306 6823
rect 11774 6538 11802 6543
rect 11662 6537 11802 6538
rect 11662 6511 11775 6537
rect 11801 6511 11802 6537
rect 11662 6510 11802 6511
rect 11774 6505 11802 6510
rect 11438 6455 11439 6481
rect 11465 6455 11466 6481
rect 11438 6449 11466 6455
rect 10822 1751 10823 1777
rect 10849 1751 10850 1777
rect 10822 1745 10850 1751
rect 11774 1834 11802 1839
rect 11214 1666 11242 1671
rect 11102 1665 11242 1666
rect 11102 1639 11215 1665
rect 11241 1639 11242 1665
rect 11102 1638 11242 1639
rect 11102 400 11130 1638
rect 11214 1633 11242 1638
rect 11774 400 11802 1806
rect 12278 1777 12306 6790
rect 12838 6537 12866 6846
rect 12838 6511 12839 6537
rect 12865 6511 12866 6537
rect 12838 2169 12866 6511
rect 13118 6537 13146 7126
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 13118 6511 13119 6537
rect 13145 6511 13146 6537
rect 13118 6505 13146 6511
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12838 2143 12839 2169
rect 12865 2143 12866 2169
rect 12838 2137 12866 2143
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12446 2058 12474 2063
rect 12446 400 12474 2030
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 8736 0 8792 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 11088 0 11144 400
rect 11760 0 11816 400
rect 12432 0 12488 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8750 19110 8778 19138
rect 9310 19137 9338 19138
rect 9310 19111 9311 19137
rect 9311 19111 9337 19137
rect 9337 19111 9338 19137
rect 9310 19110 9338 19111
rect 8414 18718 8442 18746
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9198 18745 9226 18746
rect 9198 18719 9199 18745
rect 9199 18719 9225 18745
rect 9225 18719 9226 18745
rect 9198 18718 9226 18719
rect 10430 19110 10458 19138
rect 11046 19137 11074 19138
rect 11046 19111 11047 19137
rect 11047 19111 11073 19137
rect 11073 19111 11074 19137
rect 11046 19110 11074 19111
rect 12782 19278 12810 19306
rect 13398 19278 13426 19306
rect 11438 19110 11466 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 7462 14265 7490 14266
rect 7462 14239 7463 14265
rect 7463 14239 7489 14265
rect 7489 14239 7490 14265
rect 7462 14238 7490 14239
rect 8190 14238 8218 14266
rect 7126 14182 7154 14210
rect 2086 14126 2114 14154
rect 966 11774 994 11802
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 8246 13929 8274 13930
rect 8246 13903 8247 13929
rect 8247 13903 8273 13929
rect 8273 13903 8274 13929
rect 8246 13902 8274 13903
rect 8134 13566 8162 13594
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 6454 12390 6482 12418
rect 7462 13481 7490 13482
rect 7462 13455 7463 13481
rect 7463 13455 7489 13481
rect 7489 13455 7490 13481
rect 7462 13454 7490 13455
rect 8694 13929 8722 13930
rect 8694 13903 8695 13929
rect 8695 13903 8721 13929
rect 8721 13903 8722 13929
rect 8694 13902 8722 13903
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 8862 14209 8890 14210
rect 8862 14183 8863 14209
rect 8863 14183 8889 14209
rect 8889 14183 8890 14209
rect 8862 14182 8890 14183
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 8134 12865 8162 12866
rect 8134 12839 8135 12865
rect 8135 12839 8161 12865
rect 8161 12839 8162 12865
rect 8134 12838 8162 12839
rect 8022 12782 8050 12810
rect 7126 12390 7154 12418
rect 7910 12390 7938 12418
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 4998 12025 5026 12026
rect 4998 11999 4999 12025
rect 4999 11999 5025 12025
rect 5025 11999 5026 12025
rect 4998 11998 5026 11999
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 7966 12334 7994 12362
rect 6846 12305 6874 12306
rect 6846 12279 6847 12305
rect 6847 12279 6873 12305
rect 6873 12279 6874 12305
rect 6846 12278 6874 12279
rect 6958 11998 6986 12026
rect 6398 11969 6426 11970
rect 6398 11943 6399 11969
rect 6399 11943 6425 11969
rect 6425 11943 6426 11969
rect 6398 11942 6426 11943
rect 6734 11942 6762 11970
rect 6286 11577 6314 11578
rect 6286 11551 6287 11577
rect 6287 11551 6313 11577
rect 6313 11551 6314 11577
rect 6286 11550 6314 11551
rect 2086 11494 2114 11522
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6342 11129 6370 11130
rect 6342 11103 6343 11129
rect 6343 11103 6369 11129
rect 6369 11103 6370 11129
rect 6342 11102 6370 11103
rect 5558 10793 5586 10794
rect 5558 10767 5559 10793
rect 5559 10767 5585 10793
rect 5585 10767 5586 10793
rect 5558 10766 5586 10767
rect 6846 11662 6874 11690
rect 6790 11129 6818 11130
rect 6790 11103 6791 11129
rect 6791 11103 6817 11129
rect 6817 11103 6818 11129
rect 6790 11102 6818 11103
rect 6790 10766 6818 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 7854 11998 7882 12026
rect 7182 11689 7210 11690
rect 7182 11663 7183 11689
rect 7183 11663 7209 11689
rect 7209 11663 7210 11689
rect 7182 11662 7210 11663
rect 7070 11633 7098 11634
rect 7070 11607 7071 11633
rect 7071 11607 7097 11633
rect 7097 11607 7098 11633
rect 7070 11606 7098 11607
rect 7014 11577 7042 11578
rect 7014 11551 7015 11577
rect 7015 11551 7041 11577
rect 7041 11551 7042 11577
rect 7014 11550 7042 11551
rect 7238 11606 7266 11634
rect 6958 11185 6986 11186
rect 6958 11159 6959 11185
rect 6959 11159 6985 11185
rect 6985 11159 6986 11185
rect 6958 11158 6986 11159
rect 7350 11633 7378 11634
rect 7350 11607 7351 11633
rect 7351 11607 7377 11633
rect 7377 11607 7378 11633
rect 7350 11606 7378 11607
rect 7798 11857 7826 11858
rect 7798 11831 7799 11857
rect 7799 11831 7825 11857
rect 7825 11831 7826 11857
rect 7798 11830 7826 11831
rect 7686 11606 7714 11634
rect 7294 10990 7322 11018
rect 7854 10934 7882 10962
rect 7182 10793 7210 10794
rect 7182 10767 7183 10793
rect 7183 10767 7209 10793
rect 7209 10767 7210 10793
rect 7182 10766 7210 10767
rect 7462 10766 7490 10794
rect 8190 12753 8218 12754
rect 8190 12727 8191 12753
rect 8191 12727 8217 12753
rect 8217 12727 8218 12753
rect 8190 12726 8218 12727
rect 8078 11942 8106 11970
rect 8302 12614 8330 12642
rect 8358 12446 8386 12474
rect 8246 12278 8274 12306
rect 8190 12025 8218 12026
rect 8190 11999 8191 12025
rect 8191 11999 8217 12025
rect 8217 11999 8218 12025
rect 8190 11998 8218 11999
rect 8806 13566 8834 13594
rect 8694 13510 8722 13538
rect 10710 14321 10738 14322
rect 10710 14295 10711 14321
rect 10711 14295 10737 14321
rect 10737 14295 10738 14321
rect 10710 14294 10738 14295
rect 11438 14238 11466 14266
rect 9590 13566 9618 13594
rect 8750 13481 8778 13482
rect 8750 13455 8751 13481
rect 8751 13455 8777 13481
rect 8777 13455 8778 13481
rect 8750 13454 8778 13455
rect 9478 13537 9506 13538
rect 9478 13511 9479 13537
rect 9479 13511 9505 13537
rect 9505 13511 9506 13537
rect 9478 13510 9506 13511
rect 8806 12838 8834 12866
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9030 12809 9058 12810
rect 9030 12783 9031 12809
rect 9031 12783 9057 12809
rect 9057 12783 9058 12809
rect 9030 12782 9058 12783
rect 8974 12726 9002 12754
rect 8918 12697 8946 12698
rect 8918 12671 8919 12697
rect 8919 12671 8945 12697
rect 8945 12671 8946 12697
rect 8918 12670 8946 12671
rect 8526 12334 8554 12362
rect 8750 12446 8778 12474
rect 8974 12641 9002 12642
rect 8974 12615 8975 12641
rect 8975 12615 9001 12641
rect 9001 12615 9002 12641
rect 8974 12614 9002 12615
rect 8246 11886 8274 11914
rect 8302 11774 8330 11802
rect 8134 11606 8162 11634
rect 8302 11577 8330 11578
rect 8302 11551 8303 11577
rect 8303 11551 8329 11577
rect 8329 11551 8330 11577
rect 8302 11550 8330 11551
rect 8414 11438 8442 11466
rect 8414 11185 8442 11186
rect 8414 11159 8415 11185
rect 8415 11159 8441 11185
rect 8441 11159 8442 11185
rect 8414 11158 8442 11159
rect 8750 11998 8778 12026
rect 8526 11969 8554 11970
rect 8526 11943 8527 11969
rect 8527 11943 8553 11969
rect 8553 11943 8554 11969
rect 8526 11942 8554 11943
rect 8582 11830 8610 11858
rect 8582 11662 8610 11690
rect 8638 11774 8666 11802
rect 8302 10934 8330 10962
rect 7462 10430 7490 10458
rect 7126 10206 7154 10234
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6118 9478 6146 9506
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 5726 8806 5754 8834
rect 7238 9926 7266 9954
rect 7406 10009 7434 10010
rect 7406 9983 7407 10009
rect 7407 9983 7433 10009
rect 7433 9983 7434 10009
rect 7406 9982 7434 9983
rect 7574 10289 7602 10290
rect 7574 10263 7575 10289
rect 7575 10263 7601 10289
rect 7601 10263 7602 10289
rect 7574 10262 7602 10263
rect 7854 10457 7882 10458
rect 7854 10431 7855 10457
rect 7855 10431 7881 10457
rect 7881 10431 7882 10457
rect 7854 10430 7882 10431
rect 7630 10206 7658 10234
rect 7910 10009 7938 10010
rect 7910 9983 7911 10009
rect 7911 9983 7937 10009
rect 7937 9983 7938 10009
rect 7910 9982 7938 9983
rect 7630 9953 7658 9954
rect 7630 9927 7631 9953
rect 7631 9927 7657 9953
rect 7657 9927 7658 9953
rect 7630 9926 7658 9927
rect 8470 10822 8498 10850
rect 8246 9982 8274 10010
rect 8190 9702 8218 9730
rect 8358 9982 8386 10010
rect 8358 9673 8386 9674
rect 8358 9647 8359 9673
rect 8359 9647 8385 9673
rect 8385 9647 8386 9673
rect 8358 9646 8386 9647
rect 8694 11606 8722 11634
rect 8918 11942 8946 11970
rect 8974 12278 9002 12306
rect 9422 12305 9450 12306
rect 9422 12279 9423 12305
rect 9423 12279 9449 12305
rect 9449 12279 9450 12305
rect 9422 12278 9450 12279
rect 9926 12641 9954 12642
rect 9926 12615 9927 12641
rect 9927 12615 9953 12641
rect 9953 12615 9954 12641
rect 9926 12614 9954 12615
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9646 12361 9674 12362
rect 9646 12335 9647 12361
rect 9647 12335 9673 12361
rect 9673 12335 9674 12361
rect 9646 12334 9674 12335
rect 8918 11774 8946 11802
rect 8862 11550 8890 11578
rect 8806 11521 8834 11522
rect 8806 11495 8807 11521
rect 8807 11495 8833 11521
rect 8833 11495 8834 11521
rect 8806 11494 8834 11495
rect 8918 10849 8946 10850
rect 8918 10823 8919 10849
rect 8919 10823 8945 10849
rect 8945 10823 8946 10849
rect 8918 10822 8946 10823
rect 8806 9702 8834 9730
rect 8470 9310 8498 9338
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 6790 8638 6818 8666
rect 7182 8582 7210 8610
rect 5838 8414 5866 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 966 8078 994 8106
rect 2142 8049 2170 8050
rect 2142 8023 2143 8049
rect 2143 8023 2169 8049
rect 2169 8023 2170 8049
rect 2142 8022 2170 8023
rect 1022 7742 1050 7770
rect 6902 8358 6930 8386
rect 5894 8022 5922 8050
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 6958 7910 6986 7938
rect 7350 8806 7378 8834
rect 7966 8862 7994 8890
rect 7462 8721 7490 8722
rect 7462 8695 7463 8721
rect 7463 8695 7489 8721
rect 7489 8695 7490 8721
rect 7462 8694 7490 8695
rect 7406 8582 7434 8610
rect 7406 8497 7434 8498
rect 7406 8471 7407 8497
rect 7407 8471 7433 8497
rect 7433 8471 7434 8497
rect 7406 8470 7434 8471
rect 7518 8441 7546 8442
rect 7518 8415 7519 8441
rect 7519 8415 7545 8441
rect 7545 8415 7546 8441
rect 7518 8414 7546 8415
rect 7854 8833 7882 8834
rect 7854 8807 7855 8833
rect 7855 8807 7881 8833
rect 7881 8807 7882 8833
rect 7854 8806 7882 8807
rect 7742 8721 7770 8722
rect 7742 8695 7743 8721
rect 7743 8695 7769 8721
rect 7769 8695 7770 8721
rect 7742 8694 7770 8695
rect 7798 8638 7826 8666
rect 8638 9590 8666 9618
rect 8918 9590 8946 9618
rect 9142 11270 9170 11298
rect 9142 10990 9170 11018
rect 9086 9870 9114 9898
rect 9142 10262 9170 10290
rect 8974 9646 9002 9674
rect 8750 9505 8778 9506
rect 8750 9479 8751 9505
rect 8751 9479 8777 9505
rect 8777 9479 8778 9505
rect 8750 9478 8778 9479
rect 8470 8806 8498 8834
rect 9142 9673 9170 9674
rect 9142 9647 9143 9673
rect 9143 9647 9169 9673
rect 9169 9647 9170 9673
rect 9142 9646 9170 9647
rect 9086 9590 9114 9618
rect 8918 8806 8946 8834
rect 8246 8582 8274 8610
rect 7350 8022 7378 8050
rect 7798 8441 7826 8442
rect 7798 8415 7799 8441
rect 7799 8415 7825 8441
rect 7825 8415 7826 8441
rect 7798 8414 7826 8415
rect 7910 8441 7938 8442
rect 7910 8415 7911 8441
rect 7911 8415 7937 8441
rect 7937 8415 7938 8441
rect 7910 8414 7938 8415
rect 7854 8385 7882 8386
rect 7854 8359 7855 8385
rect 7855 8359 7881 8385
rect 7881 8359 7882 8385
rect 7854 8358 7882 8359
rect 7742 8302 7770 8330
rect 7798 8078 7826 8106
rect 9254 10038 9282 10066
rect 9366 10009 9394 10010
rect 9366 9983 9367 10009
rect 9367 9983 9393 10009
rect 9393 9983 9394 10009
rect 9366 9982 9394 9983
rect 9310 9870 9338 9898
rect 9814 11913 9842 11914
rect 9814 11887 9815 11913
rect 9815 11887 9841 11913
rect 9841 11887 9842 11913
rect 9814 11886 9842 11887
rect 9590 11494 9618 11522
rect 9478 10206 9506 10234
rect 9646 10038 9674 10066
rect 9254 8889 9282 8890
rect 9254 8863 9255 8889
rect 9255 8863 9281 8889
rect 9281 8863 9282 8889
rect 9254 8862 9282 8863
rect 9422 9534 9450 9562
rect 9702 9926 9730 9954
rect 11270 13985 11298 13986
rect 11270 13959 11271 13985
rect 11271 13959 11297 13985
rect 11297 13959 11298 13985
rect 11270 13958 11298 13959
rect 10822 13929 10850 13930
rect 10822 13903 10823 13929
rect 10823 13903 10849 13929
rect 10849 13903 10850 13929
rect 10822 13902 10850 13903
rect 11214 13929 11242 13930
rect 11214 13903 11215 13929
rect 11215 13903 11241 13929
rect 11241 13903 11242 13929
rect 11214 13902 11242 13903
rect 10878 13566 10906 13594
rect 12334 14321 12362 14322
rect 12334 14295 12335 14321
rect 12335 14295 12361 14321
rect 12361 14295 12362 14321
rect 12334 14294 12362 14295
rect 12110 13958 12138 13986
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 20118 17150 20146 17178
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 11046 13286 11074 13314
rect 11438 13286 11466 13314
rect 12726 13286 12754 13314
rect 10654 12697 10682 12698
rect 10654 12671 10655 12697
rect 10655 12671 10681 12697
rect 10681 12671 10682 12697
rect 10654 12670 10682 12671
rect 10262 12417 10290 12418
rect 10262 12391 10263 12417
rect 10263 12391 10289 12417
rect 10289 12391 10290 12417
rect 10262 12390 10290 12391
rect 10150 12361 10178 12362
rect 10150 12335 10151 12361
rect 10151 12335 10177 12361
rect 10177 12335 10178 12361
rect 10150 12334 10178 12335
rect 10710 12166 10738 12194
rect 10822 12278 10850 12306
rect 10150 11998 10178 12026
rect 10654 12025 10682 12026
rect 10654 11999 10655 12025
rect 10655 11999 10681 12025
rect 10681 11999 10682 12025
rect 10654 11998 10682 11999
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10374 11857 10402 11858
rect 10374 11831 10375 11857
rect 10375 11831 10401 11857
rect 10401 11831 10402 11857
rect 10374 11830 10402 11831
rect 10262 11662 10290 11690
rect 10262 11214 10290 11242
rect 10206 11158 10234 11186
rect 9926 11073 9954 11074
rect 9926 11047 9927 11073
rect 9927 11047 9953 11073
rect 9953 11047 9954 11073
rect 9926 11046 9954 11047
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10206 10934 10234 10962
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9982 10038 10010 10066
rect 10710 11129 10738 11130
rect 10710 11103 10711 11129
rect 10711 11103 10737 11129
rect 10737 11103 10738 11129
rect 10710 11102 10738 11103
rect 10262 9982 10290 10010
rect 9534 9310 9562 9338
rect 9646 9422 9674 9450
rect 9422 9086 9450 9114
rect 8862 8078 8890 8106
rect 7574 7937 7602 7938
rect 7574 7911 7575 7937
rect 7575 7911 7601 7937
rect 7601 7911 7602 7937
rect 7574 7910 7602 7911
rect 7742 7574 7770 7602
rect 7574 7126 7602 7154
rect 8806 7713 8834 7714
rect 8806 7687 8807 7713
rect 8807 7687 8833 7713
rect 8833 7687 8834 7713
rect 8806 7686 8834 7687
rect 9254 8358 9282 8386
rect 8862 7601 8890 7602
rect 8862 7575 8863 7601
rect 8863 7575 8889 7601
rect 8889 7575 8890 7601
rect 8862 7574 8890 7575
rect 9030 7462 9058 7490
rect 9198 7462 9226 7490
rect 8750 7126 8778 7154
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 9254 7209 9282 7210
rect 9254 7183 9255 7209
rect 9255 7183 9281 7209
rect 9281 7183 9282 7209
rect 9254 7182 9282 7183
rect 9870 9702 9898 9730
rect 9870 9478 9898 9506
rect 10654 11046 10682 11074
rect 10710 10934 10738 10962
rect 11102 12166 11130 12194
rect 11046 11969 11074 11970
rect 11046 11943 11047 11969
rect 11047 11943 11073 11969
rect 11073 11943 11074 11969
rect 11046 11942 11074 11943
rect 10878 11073 10906 11074
rect 10878 11047 10879 11073
rect 10879 11047 10905 11073
rect 10905 11047 10906 11073
rect 10878 11046 10906 11047
rect 11158 11689 11186 11690
rect 11158 11663 11159 11689
rect 11159 11663 11185 11689
rect 11185 11663 11186 11689
rect 11158 11662 11186 11663
rect 11214 11830 11242 11858
rect 11102 11270 11130 11298
rect 11046 11046 11074 11074
rect 10822 10710 10850 10738
rect 10430 9926 10458 9954
rect 10374 9646 10402 9674
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10150 9198 10178 9226
rect 10318 9478 10346 9506
rect 10710 9617 10738 9618
rect 10710 9591 10711 9617
rect 10711 9591 10737 9617
rect 10737 9591 10738 9617
rect 10710 9590 10738 9591
rect 10486 9281 10514 9282
rect 10486 9255 10487 9281
rect 10487 9255 10513 9281
rect 10513 9255 10514 9281
rect 10486 9254 10514 9255
rect 10654 9310 10682 9338
rect 10878 10094 10906 10122
rect 10934 9702 10962 9730
rect 11326 12390 11354 12418
rect 11438 12614 11466 12642
rect 11382 11942 11410 11970
rect 11382 11774 11410 11802
rect 11438 11718 11466 11746
rect 11494 11830 11522 11858
rect 11438 11550 11466 11578
rect 11662 13145 11690 13146
rect 11662 13119 11663 13145
rect 11663 13119 11689 13145
rect 11689 13119 11690 13145
rect 11662 13118 11690 13119
rect 12614 13145 12642 13146
rect 12614 13119 12615 13145
rect 12615 13119 12641 13145
rect 12641 13119 12642 13145
rect 12614 13118 12642 13119
rect 11662 12473 11690 12474
rect 11662 12447 11663 12473
rect 11663 12447 11689 12473
rect 11689 12447 11690 12473
rect 11662 12446 11690 12447
rect 12110 12473 12138 12474
rect 12110 12447 12111 12473
rect 12111 12447 12137 12473
rect 12137 12447 12138 12473
rect 12110 12446 12138 12447
rect 13118 13286 13146 13314
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 12446 12446 12474 12474
rect 11550 11774 11578 11802
rect 11662 11718 11690 11746
rect 11382 11241 11410 11242
rect 11382 11215 11383 11241
rect 11383 11215 11409 11241
rect 11409 11215 11410 11241
rect 11382 11214 11410 11215
rect 11214 11158 11242 11186
rect 11158 10401 11186 10402
rect 11158 10375 11159 10401
rect 11159 10375 11185 10401
rect 11185 10375 11186 10401
rect 11158 10374 11186 10375
rect 11102 9534 11130 9562
rect 10990 9478 11018 9506
rect 11158 9478 11186 9506
rect 11102 9254 11130 9282
rect 10934 9225 10962 9226
rect 10934 9199 10935 9225
rect 10935 9199 10961 9225
rect 10961 9199 10962 9225
rect 10934 9198 10962 9199
rect 10766 8918 10794 8946
rect 10822 8833 10850 8834
rect 10822 8807 10823 8833
rect 10823 8807 10849 8833
rect 10849 8807 10850 8833
rect 10822 8806 10850 8807
rect 9646 7350 9674 7378
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10654 8553 10682 8554
rect 10654 8527 10655 8553
rect 10655 8527 10681 8553
rect 10681 8527 10682 8553
rect 10654 8526 10682 8527
rect 10878 8414 10906 8442
rect 10710 7910 10738 7938
rect 10822 7966 10850 7994
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9926 7601 9954 7602
rect 9926 7575 9927 7601
rect 9927 7575 9953 7601
rect 9953 7575 9954 7601
rect 9926 7574 9954 7575
rect 10822 7574 10850 7602
rect 9982 7377 10010 7378
rect 9982 7351 9983 7377
rect 9983 7351 10009 7377
rect 10009 7351 10010 7377
rect 9982 7350 10010 7351
rect 9814 7294 9842 7322
rect 9758 7265 9786 7266
rect 9758 7239 9759 7265
rect 9759 7239 9785 7265
rect 9785 7239 9786 7265
rect 9758 7238 9786 7239
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9814 6790 9842 6818
rect 9310 6734 9338 6762
rect 8750 2030 8778 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9254 2057 9282 2058
rect 9254 2031 9255 2057
rect 9255 2031 9281 2057
rect 9281 2031 9282 2057
rect 9254 2030 9282 2031
rect 10430 7294 10458 7322
rect 10374 7153 10402 7154
rect 10374 7127 10375 7153
rect 10375 7127 10401 7153
rect 10401 7127 10402 7153
rect 10374 7126 10402 7127
rect 10542 7182 10570 7210
rect 10150 6817 10178 6818
rect 10150 6791 10151 6817
rect 10151 6791 10177 6817
rect 10177 6791 10178 6817
rect 10150 6790 10178 6791
rect 10598 6761 10626 6762
rect 10598 6735 10599 6761
rect 10599 6735 10625 6761
rect 10625 6735 10626 6761
rect 10598 6734 10626 6735
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10094 2030 10122 2058
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 10710 2057 10738 2058
rect 10710 2031 10711 2057
rect 10711 2031 10737 2057
rect 10737 2031 10738 2057
rect 10710 2030 10738 2031
rect 11326 10934 11354 10962
rect 11382 10094 11410 10122
rect 11830 11662 11858 11690
rect 11718 11214 11746 11242
rect 11886 11633 11914 11634
rect 11886 11607 11887 11633
rect 11887 11607 11913 11633
rect 11913 11607 11914 11633
rect 11886 11606 11914 11607
rect 12110 11886 12138 11914
rect 12390 11830 12418 11858
rect 11662 11102 11690 11130
rect 11942 10990 11970 11018
rect 12166 11046 12194 11074
rect 11606 10654 11634 10682
rect 12110 10038 12138 10066
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 12894 11913 12922 11914
rect 12894 11887 12895 11913
rect 12895 11887 12921 11913
rect 12921 11887 12922 11913
rect 12894 11886 12922 11887
rect 12278 11521 12306 11522
rect 12278 11495 12279 11521
rect 12279 11495 12305 11521
rect 12305 11495 12306 11521
rect 12278 11494 12306 11495
rect 12838 11326 12866 11354
rect 12502 11214 12530 11242
rect 12278 11185 12306 11186
rect 12278 11159 12279 11185
rect 12279 11159 12305 11185
rect 12305 11159 12306 11185
rect 12278 11158 12306 11159
rect 11438 9702 11466 9730
rect 11326 9617 11354 9618
rect 11326 9591 11327 9617
rect 11327 9591 11353 9617
rect 11353 9591 11354 9617
rect 11326 9590 11354 9591
rect 11046 7966 11074 7994
rect 11214 8526 11242 8554
rect 10990 7910 11018 7938
rect 11046 7321 11074 7322
rect 11046 7295 11047 7321
rect 11047 7295 11073 7321
rect 11073 7295 11074 7321
rect 11046 7294 11074 7295
rect 11382 9310 11410 9338
rect 11438 9254 11466 9282
rect 11718 9673 11746 9674
rect 11718 9647 11719 9673
rect 11719 9647 11745 9673
rect 11745 9647 11746 9673
rect 11718 9646 11746 9647
rect 11662 9534 11690 9562
rect 11494 8945 11522 8946
rect 11494 8919 11495 8945
rect 11495 8919 11521 8945
rect 11521 8919 11522 8945
rect 11494 8918 11522 8919
rect 11326 8833 11354 8834
rect 11326 8807 11327 8833
rect 11327 8807 11353 8833
rect 11353 8807 11354 8833
rect 11326 8806 11354 8807
rect 11550 8526 11578 8554
rect 12390 10094 12418 10122
rect 13006 11326 13034 11354
rect 13286 11942 13314 11970
rect 13958 11969 13986 11970
rect 13958 11943 13959 11969
rect 13959 11943 13985 11969
rect 13985 11943 13986 11969
rect 13958 11942 13986 11943
rect 14294 11942 14322 11970
rect 13398 11857 13426 11858
rect 13398 11831 13399 11857
rect 13399 11831 13425 11857
rect 13425 11831 13426 11857
rect 13398 11830 13426 11831
rect 14070 11857 14098 11858
rect 14070 11831 14071 11857
rect 14071 11831 14097 11857
rect 14097 11831 14098 11857
rect 14070 11830 14098 11831
rect 13230 11521 13258 11522
rect 13230 11495 13231 11521
rect 13231 11495 13257 11521
rect 13257 11495 13258 11521
rect 13230 11494 13258 11495
rect 13006 10990 13034 11018
rect 12838 10905 12866 10906
rect 12838 10879 12839 10905
rect 12839 10879 12865 10905
rect 12865 10879 12866 10905
rect 12838 10878 12866 10879
rect 12950 10849 12978 10850
rect 12950 10823 12951 10849
rect 12951 10823 12977 10849
rect 12977 10823 12978 10849
rect 12950 10822 12978 10823
rect 12446 10038 12474 10066
rect 12446 9617 12474 9618
rect 12446 9591 12447 9617
rect 12447 9591 12473 9617
rect 12473 9591 12474 9617
rect 12446 9590 12474 9591
rect 12950 10654 12978 10682
rect 12726 10094 12754 10122
rect 13062 11102 13090 11130
rect 13902 11550 13930 11578
rect 13174 10905 13202 10906
rect 13174 10879 13175 10905
rect 13175 10879 13201 10905
rect 13201 10879 13202 10905
rect 13174 10878 13202 10879
rect 13398 10990 13426 11018
rect 13118 10737 13146 10738
rect 13118 10711 13119 10737
rect 13119 10711 13145 10737
rect 13145 10711 13146 10737
rect 13118 10710 13146 10711
rect 12614 9534 12642 9562
rect 13062 9702 13090 9730
rect 12166 9281 12194 9282
rect 12166 9255 12167 9281
rect 12167 9255 12193 9281
rect 12193 9255 12194 9281
rect 12166 9254 12194 9255
rect 11718 9198 11746 9226
rect 11998 9142 12026 9170
rect 12558 9142 12586 9170
rect 13174 9505 13202 9506
rect 13174 9479 13175 9505
rect 13175 9479 13201 9505
rect 13201 9479 13202 9505
rect 13174 9478 13202 9479
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 18830 11830 18858 11858
rect 20006 11774 20034 11802
rect 14294 11241 14322 11242
rect 14294 11215 14295 11241
rect 14295 11215 14321 11241
rect 14321 11215 14322 11241
rect 14294 11214 14322 11215
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 20006 11102 20034 11130
rect 14518 10990 14546 11018
rect 14294 10822 14322 10850
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 12670 9086 12698 9114
rect 12782 8414 12810 8442
rect 12838 9198 12866 9226
rect 12894 8918 12922 8946
rect 13118 9086 13146 9114
rect 13398 9225 13426 9226
rect 13398 9199 13399 9225
rect 13399 9199 13425 9225
rect 13425 9199 13426 9225
rect 13398 9198 13426 9199
rect 11998 8358 12026 8386
rect 13734 9561 13762 9562
rect 13734 9535 13735 9561
rect 13735 9535 13761 9561
rect 13761 9535 13762 9561
rect 13734 9534 13762 9535
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14686 9534 14714 9562
rect 14798 9590 14826 9618
rect 14854 9534 14882 9562
rect 13622 9086 13650 9114
rect 13510 8862 13538 8890
rect 13454 8777 13482 8778
rect 13454 8751 13455 8777
rect 13455 8751 13481 8777
rect 13481 8751 13482 8777
rect 13454 8750 13482 8751
rect 13398 8694 13426 8722
rect 15022 9534 15050 9562
rect 15134 9505 15162 9506
rect 15134 9479 15135 9505
rect 15135 9479 15161 9505
rect 15161 9479 15162 9505
rect 15134 9478 15162 9479
rect 20006 10094 20034 10122
rect 20006 9758 20034 9786
rect 18942 9702 18970 9730
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 18774 9478 18802 9506
rect 20006 9422 20034 9450
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14182 8862 14210 8890
rect 13790 8806 13818 8834
rect 14462 8806 14490 8834
rect 13902 8777 13930 8778
rect 13902 8751 13903 8777
rect 13903 8751 13929 8777
rect 13929 8751 13930 8777
rect 13902 8750 13930 8751
rect 14070 8721 14098 8722
rect 14070 8695 14071 8721
rect 14071 8695 14097 8721
rect 14097 8695 14098 8721
rect 14070 8694 14098 8695
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 14518 8694 14546 8722
rect 13734 8049 13762 8050
rect 13734 8023 13735 8049
rect 13735 8023 13761 8049
rect 13761 8023 13762 8049
rect 13734 8022 13762 8023
rect 14294 8022 14322 8050
rect 13230 7686 13258 7714
rect 11438 7406 11466 7434
rect 11382 7321 11410 7322
rect 11382 7295 11383 7321
rect 11383 7295 11409 7321
rect 11409 7295 11410 7321
rect 11382 7294 11410 7295
rect 11102 7238 11130 7266
rect 11270 7265 11298 7266
rect 11270 7239 11271 7265
rect 11271 7239 11297 7265
rect 11297 7239 11298 7265
rect 11270 7238 11298 7239
rect 10878 6873 10906 6874
rect 10878 6847 10879 6873
rect 10879 6847 10905 6873
rect 10905 6847 10906 6873
rect 10878 6846 10906 6847
rect 11438 7126 11466 7154
rect 11718 7406 11746 7434
rect 12614 7350 12642 7378
rect 11606 7126 11634 7154
rect 11438 6846 11466 6874
rect 11046 6790 11074 6818
rect 11942 7265 11970 7266
rect 11942 7239 11943 7265
rect 11943 7239 11969 7265
rect 11969 7239 11970 7265
rect 11942 7238 11970 7239
rect 11718 7182 11746 7210
rect 12390 7153 12418 7154
rect 12390 7127 12391 7153
rect 12391 7127 12417 7153
rect 12417 7127 12418 7153
rect 12390 7126 12418 7127
rect 12670 7238 12698 7266
rect 13174 7350 13202 7378
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 18830 8049 18858 8050
rect 18830 8023 18831 8049
rect 18831 8023 18857 8049
rect 18857 8023 18858 8049
rect 18830 8022 18858 8023
rect 20006 7742 20034 7770
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 12838 7126 12866 7154
rect 13118 7126 13146 7154
rect 12278 6817 12306 6818
rect 12278 6791 12279 6817
rect 12279 6791 12305 6817
rect 12305 6791 12306 6817
rect 12278 6790 12306 6791
rect 11774 1806 11802 1834
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12446 2030 12474 2058
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 12777 19278 12782 19306
rect 12810 19278 13398 19306
rect 13426 19278 13431 19306
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8745 19110 8750 19138
rect 8778 19110 9310 19138
rect 9338 19110 9343 19138
rect 10425 19110 10430 19138
rect 10458 19110 11046 19138
rect 11074 19110 11079 19138
rect 11433 19110 11438 19138
rect 11466 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8409 18718 8414 18746
rect 8442 18718 9198 18746
rect 9226 18718 9231 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 20600 17178 21000 17192
rect 20113 17150 20118 17178
rect 20146 17150 21000 17178
rect 20600 17136 21000 17150
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 10705 14294 10710 14322
rect 10738 14294 12334 14322
rect 12362 14294 12367 14322
rect 11438 14266 11466 14294
rect 7457 14238 7462 14266
rect 7490 14238 8190 14266
rect 8218 14238 8223 14266
rect 11433 14238 11438 14266
rect 11466 14238 11471 14266
rect 7121 14182 7126 14210
rect 7154 14182 8862 14210
rect 8890 14182 8895 14210
rect 0 14154 400 14168
rect 0 14126 2086 14154
rect 2114 14126 2119 14154
rect 0 14112 400 14126
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 11265 13958 11270 13986
rect 11298 13958 12110 13986
rect 12138 13958 12143 13986
rect 8241 13902 8246 13930
rect 8274 13902 8694 13930
rect 8722 13902 8727 13930
rect 10817 13902 10822 13930
rect 10850 13902 11214 13930
rect 11242 13902 11247 13930
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 8129 13566 8134 13594
rect 8162 13566 8806 13594
rect 8834 13566 9590 13594
rect 9618 13566 10878 13594
rect 10906 13566 10911 13594
rect 8689 13510 8694 13538
rect 8722 13510 9478 13538
rect 9506 13510 9511 13538
rect 7457 13454 7462 13482
rect 7490 13454 8750 13482
rect 8778 13454 8783 13482
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 11041 13286 11046 13314
rect 11074 13286 11438 13314
rect 11466 13286 12726 13314
rect 12754 13286 13118 13314
rect 13146 13286 13151 13314
rect 11657 13118 11662 13146
rect 11690 13118 12614 13146
rect 12642 13118 12647 13146
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 8129 12838 8134 12866
rect 8162 12838 8806 12866
rect 8834 12838 8839 12866
rect 8017 12782 8022 12810
rect 8050 12782 9030 12810
rect 9058 12782 9063 12810
rect 8185 12726 8190 12754
rect 8218 12726 8974 12754
rect 9002 12726 9007 12754
rect 8913 12670 8918 12698
rect 8946 12670 10654 12698
rect 10682 12670 10687 12698
rect 8297 12614 8302 12642
rect 8330 12614 8974 12642
rect 9002 12614 9007 12642
rect 9921 12614 9926 12642
rect 9954 12614 11438 12642
rect 11466 12614 11471 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 8353 12446 8358 12474
rect 8386 12446 8750 12474
rect 8778 12446 8783 12474
rect 11657 12446 11662 12474
rect 11690 12446 12110 12474
rect 12138 12446 12446 12474
rect 12474 12446 12479 12474
rect 6449 12390 6454 12418
rect 6482 12390 7126 12418
rect 7154 12390 7910 12418
rect 7938 12390 7943 12418
rect 10257 12390 10262 12418
rect 10290 12390 11326 12418
rect 11354 12390 11359 12418
rect 7961 12334 7966 12362
rect 7994 12334 8526 12362
rect 8554 12334 9646 12362
rect 9674 12334 10150 12362
rect 10178 12334 10183 12362
rect 6841 12278 6846 12306
rect 6874 12278 8246 12306
rect 8274 12278 8279 12306
rect 8969 12278 8974 12306
rect 9002 12278 9422 12306
rect 9450 12278 10822 12306
rect 10850 12278 10855 12306
rect 10705 12166 10710 12194
rect 10738 12166 11102 12194
rect 11130 12166 11135 12194
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 4186 11998 4998 12026
rect 5026 11998 6958 12026
rect 6986 11998 6991 12026
rect 7849 11998 7854 12026
rect 7882 11998 8190 12026
rect 8218 11998 8750 12026
rect 8778 11998 8783 12026
rect 10145 11998 10150 12026
rect 10178 11998 10654 12026
rect 10682 11998 10687 12026
rect 4186 11970 4214 11998
rect 2137 11942 2142 11970
rect 2170 11942 4214 11970
rect 6393 11942 6398 11970
rect 6426 11942 6734 11970
rect 6762 11942 6767 11970
rect 8073 11942 8078 11970
rect 8106 11942 8526 11970
rect 8554 11942 8559 11970
rect 8913 11942 8918 11970
rect 8946 11942 11046 11970
rect 11074 11942 11382 11970
rect 11410 11942 11415 11970
rect 13281 11942 13286 11970
rect 13314 11942 13958 11970
rect 13986 11942 14294 11970
rect 14322 11942 18830 11970
rect 18858 11942 18863 11970
rect 8241 11886 8246 11914
rect 8274 11886 9814 11914
rect 9842 11886 9847 11914
rect 12105 11886 12110 11914
rect 12138 11886 12894 11914
rect 12922 11886 12927 11914
rect 7793 11830 7798 11858
rect 7826 11830 8582 11858
rect 8610 11830 8615 11858
rect 10369 11830 10374 11858
rect 10402 11830 11214 11858
rect 11242 11830 11494 11858
rect 11522 11830 11527 11858
rect 12385 11830 12390 11858
rect 12418 11830 13398 11858
rect 13426 11830 13431 11858
rect 14065 11830 14070 11858
rect 14098 11830 18830 11858
rect 18858 11830 18863 11858
rect 0 11802 400 11816
rect 20600 11802 21000 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 8297 11774 8302 11802
rect 8330 11774 8638 11802
rect 8666 11774 8918 11802
rect 8946 11774 8951 11802
rect 11377 11774 11382 11802
rect 11410 11774 11550 11802
rect 11578 11774 11583 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 11433 11718 11438 11746
rect 11466 11718 11662 11746
rect 11690 11718 11695 11746
rect 6841 11662 6846 11690
rect 6874 11662 7182 11690
rect 7210 11662 7215 11690
rect 8577 11662 8582 11690
rect 8610 11662 10262 11690
rect 10290 11662 10295 11690
rect 11153 11662 11158 11690
rect 11186 11662 11830 11690
rect 11858 11662 11863 11690
rect 10262 11634 10290 11662
rect 7065 11606 7070 11634
rect 7098 11606 7238 11634
rect 7266 11606 7271 11634
rect 7345 11606 7350 11634
rect 7378 11606 7686 11634
rect 7714 11606 8134 11634
rect 8162 11606 8694 11634
rect 8722 11606 8727 11634
rect 10262 11606 11886 11634
rect 11914 11606 11919 11634
rect 6281 11550 6286 11578
rect 6314 11550 7014 11578
rect 7042 11550 7047 11578
rect 8297 11550 8302 11578
rect 8330 11550 8862 11578
rect 8890 11550 8895 11578
rect 11433 11550 11438 11578
rect 11466 11550 13902 11578
rect 13930 11550 13935 11578
rect 2081 11494 2086 11522
rect 2114 11494 8806 11522
rect 8834 11494 9590 11522
rect 9618 11494 9623 11522
rect 11438 11466 11466 11550
rect 12273 11494 12278 11522
rect 12306 11494 13230 11522
rect 13258 11494 13263 11522
rect 20600 11466 21000 11480
rect 8409 11438 8414 11466
rect 8442 11438 11466 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 12833 11326 12838 11354
rect 12866 11326 13006 11354
rect 13034 11326 13039 11354
rect 9137 11270 9142 11298
rect 9170 11270 11102 11298
rect 11130 11270 11135 11298
rect 10257 11214 10262 11242
rect 10290 11214 11382 11242
rect 11410 11214 11415 11242
rect 11713 11214 11718 11242
rect 11746 11214 12502 11242
rect 12530 11214 12535 11242
rect 14289 11214 14294 11242
rect 14322 11214 15974 11242
rect 15946 11186 15974 11214
rect 6953 11158 6958 11186
rect 6986 11158 8414 11186
rect 8442 11158 8447 11186
rect 10201 11158 10206 11186
rect 10234 11158 11214 11186
rect 11242 11158 12278 11186
rect 12306 11158 12311 11186
rect 15946 11158 18830 11186
rect 18858 11158 18863 11186
rect 20600 11130 21000 11144
rect 6337 11102 6342 11130
rect 6370 11102 6790 11130
rect 6818 11102 6823 11130
rect 10705 11102 10710 11130
rect 10738 11102 11662 11130
rect 11690 11102 13062 11130
rect 13090 11102 13095 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 9921 11046 9926 11074
rect 9954 11046 10654 11074
rect 10682 11046 10687 11074
rect 10873 11046 10878 11074
rect 10906 11046 11046 11074
rect 11074 11046 12166 11074
rect 12194 11046 12199 11074
rect 10654 11018 10682 11046
rect 7289 10990 7294 11018
rect 7322 10990 9142 11018
rect 9170 10990 9175 11018
rect 10654 10990 11942 11018
rect 11970 10990 11975 11018
rect 13001 10990 13006 11018
rect 13034 10990 13398 11018
rect 13426 10990 14518 11018
rect 14546 10990 14551 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7849 10934 7854 10962
rect 7882 10934 8302 10962
rect 8330 10934 8335 10962
rect 10201 10934 10206 10962
rect 10234 10934 10710 10962
rect 10738 10934 11326 10962
rect 11354 10934 11359 10962
rect 12833 10878 12838 10906
rect 12866 10878 13174 10906
rect 13202 10878 13207 10906
rect 8465 10822 8470 10850
rect 8498 10822 8918 10850
rect 8946 10822 8951 10850
rect 12945 10822 12950 10850
rect 12978 10822 14294 10850
rect 14322 10822 14327 10850
rect 5553 10766 5558 10794
rect 5586 10766 6790 10794
rect 6818 10766 7182 10794
rect 7210 10766 7462 10794
rect 7490 10766 7495 10794
rect 10817 10710 10822 10738
rect 10850 10710 13118 10738
rect 13146 10710 13151 10738
rect 11601 10654 11606 10682
rect 11634 10654 12950 10682
rect 12978 10654 12983 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7457 10430 7462 10458
rect 7490 10430 7854 10458
rect 7882 10430 7887 10458
rect 10033 10374 10038 10402
rect 10066 10374 11158 10402
rect 11186 10374 11191 10402
rect 7569 10262 7574 10290
rect 7602 10262 9142 10290
rect 9170 10262 9175 10290
rect 7121 10206 7126 10234
rect 7154 10206 7630 10234
rect 7658 10206 9478 10234
rect 9506 10206 9511 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 20600 10122 21000 10136
rect 10873 10094 10878 10122
rect 10906 10094 11382 10122
rect 11410 10094 11415 10122
rect 12385 10094 12390 10122
rect 12418 10094 12726 10122
rect 12754 10094 12759 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 20600 10080 21000 10094
rect 9249 10038 9254 10066
rect 9282 10038 9646 10066
rect 9674 10038 9982 10066
rect 10010 10038 12110 10066
rect 12138 10038 12446 10066
rect 12474 10038 12479 10066
rect 7401 9982 7406 10010
rect 7434 9982 7910 10010
rect 7938 9982 8246 10010
rect 8274 9982 8279 10010
rect 8353 9982 8358 10010
rect 8386 9982 9366 10010
rect 9394 9982 10262 10010
rect 10290 9982 10295 10010
rect 7233 9926 7238 9954
rect 7266 9926 7630 9954
rect 7658 9926 9702 9954
rect 9730 9926 10430 9954
rect 10458 9926 10463 9954
rect 9081 9870 9086 9898
rect 9114 9870 9310 9898
rect 9338 9870 9343 9898
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 8185 9702 8190 9730
rect 8218 9702 8806 9730
rect 8834 9702 9870 9730
rect 9898 9702 9903 9730
rect 10929 9702 10934 9730
rect 10962 9702 11438 9730
rect 11466 9702 13062 9730
rect 13090 9702 13095 9730
rect 15946 9702 18942 9730
rect 18970 9702 18975 9730
rect 8353 9646 8358 9674
rect 8386 9646 8974 9674
rect 9002 9646 9007 9674
rect 9137 9646 9142 9674
rect 9170 9646 10374 9674
rect 10402 9646 11718 9674
rect 11746 9646 11751 9674
rect 15946 9618 15974 9702
rect 8633 9590 8638 9618
rect 8666 9590 8918 9618
rect 8946 9590 9086 9618
rect 9114 9590 10710 9618
rect 10738 9590 10743 9618
rect 11321 9590 11326 9618
rect 11354 9590 12446 9618
rect 12474 9590 12479 9618
rect 14793 9590 14798 9618
rect 14826 9590 15974 9618
rect 18825 9590 18830 9618
rect 18858 9590 18863 9618
rect 18830 9562 18858 9590
rect 9417 9534 9422 9562
rect 9450 9534 11102 9562
rect 11130 9534 11135 9562
rect 11657 9534 11662 9562
rect 11690 9534 12614 9562
rect 12642 9534 12647 9562
rect 13729 9534 13734 9562
rect 13762 9534 14686 9562
rect 14714 9534 14854 9562
rect 14882 9534 15022 9562
rect 15050 9534 18858 9562
rect 6113 9478 6118 9506
rect 6146 9478 8750 9506
rect 8778 9478 8783 9506
rect 9646 9478 9870 9506
rect 9898 9478 9903 9506
rect 10313 9478 10318 9506
rect 10346 9478 10990 9506
rect 11018 9478 11158 9506
rect 11186 9478 13174 9506
rect 13202 9478 13207 9506
rect 15129 9478 15134 9506
rect 15162 9478 18774 9506
rect 18802 9478 18807 9506
rect 9646 9450 9674 9478
rect 20600 9450 21000 9464
rect 9641 9422 9646 9450
rect 9674 9422 9679 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 8465 9310 8470 9338
rect 8498 9310 9534 9338
rect 9562 9310 10654 9338
rect 10682 9310 11382 9338
rect 11410 9310 11415 9338
rect 10481 9254 10486 9282
rect 10514 9254 11102 9282
rect 11130 9254 11135 9282
rect 11433 9254 11438 9282
rect 11466 9254 12166 9282
rect 12194 9254 12199 9282
rect 9422 9198 10150 9226
rect 10178 9198 10934 9226
rect 10962 9198 10967 9226
rect 11713 9198 11718 9226
rect 11746 9198 12838 9226
rect 12866 9198 13398 9226
rect 13426 9198 13431 9226
rect 15946 9198 18830 9226
rect 18858 9198 18863 9226
rect 9422 9114 9450 9198
rect 9417 9086 9422 9114
rect 9450 9086 9455 9114
rect 10934 9058 10962 9198
rect 15946 9170 15974 9198
rect 11993 9142 11998 9170
rect 12026 9142 12558 9170
rect 12586 9142 12591 9170
rect 13118 9142 15974 9170
rect 13118 9114 13146 9142
rect 20600 9114 21000 9128
rect 12665 9086 12670 9114
rect 12698 9086 13118 9114
rect 13146 9086 13151 9114
rect 13426 9086 13622 9114
rect 13650 9086 13655 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 13426 9058 13454 9086
rect 20600 9072 21000 9086
rect 10934 9030 13454 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 10761 8918 10766 8946
rect 10794 8918 11494 8946
rect 11522 8918 12894 8946
rect 12922 8918 12927 8946
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 7961 8862 7966 8890
rect 7994 8862 9254 8890
rect 9282 8862 9287 8890
rect 9366 8862 13510 8890
rect 13538 8862 14182 8890
rect 14210 8862 14215 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 9366 8834 9394 8862
rect 2137 8806 2142 8834
rect 2170 8806 5726 8834
rect 5754 8806 7350 8834
rect 7378 8806 7383 8834
rect 7849 8806 7854 8834
rect 7882 8806 8470 8834
rect 8498 8806 8503 8834
rect 8913 8806 8918 8834
rect 8946 8806 9394 8834
rect 10817 8806 10822 8834
rect 10850 8806 11326 8834
rect 11354 8806 11359 8834
rect 13785 8806 13790 8834
rect 13818 8806 14462 8834
rect 14490 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 0 8750 994 8778
rect 13449 8750 13454 8778
rect 13482 8750 13902 8778
rect 13930 8750 13935 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 0 8736 400 8750
rect 20600 8736 21000 8750
rect 7457 8694 7462 8722
rect 7490 8694 7742 8722
rect 7770 8694 7775 8722
rect 13393 8694 13398 8722
rect 13426 8694 14070 8722
rect 14098 8694 14518 8722
rect 14546 8694 14551 8722
rect 6785 8638 6790 8666
rect 6818 8638 7798 8666
rect 7826 8638 7831 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7177 8582 7182 8610
rect 7210 8582 7406 8610
rect 7434 8582 8246 8610
rect 8274 8582 8279 8610
rect 10649 8526 10654 8554
rect 10682 8526 11214 8554
rect 11242 8526 11550 8554
rect 11578 8526 11583 8554
rect 5838 8470 7406 8498
rect 7434 8470 7439 8498
rect 5838 8442 5866 8470
rect 2137 8414 2142 8442
rect 2170 8414 5838 8442
rect 5866 8414 5871 8442
rect 7513 8414 7518 8442
rect 7546 8414 7798 8442
rect 7826 8414 7831 8442
rect 7905 8414 7910 8442
rect 7938 8414 10878 8442
rect 10906 8414 12782 8442
rect 12810 8414 12815 8442
rect 6897 8358 6902 8386
rect 6930 8358 7854 8386
rect 7882 8358 7887 8386
rect 9249 8358 9254 8386
rect 9282 8358 11998 8386
rect 12026 8358 12031 8386
rect 9254 8330 9282 8358
rect 7737 8302 7742 8330
rect 7770 8302 9282 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 0 8106 400 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 7793 8078 7798 8106
rect 7826 8078 8862 8106
rect 8890 8078 8895 8106
rect 0 8064 400 8078
rect 2137 8022 2142 8050
rect 2170 8022 5894 8050
rect 5922 8022 7350 8050
rect 7378 8022 7383 8050
rect 13729 8022 13734 8050
rect 13762 8022 14294 8050
rect 14322 8022 18830 8050
rect 18858 8022 18863 8050
rect 10817 7966 10822 7994
rect 10850 7966 11046 7994
rect 11074 7966 11079 7994
rect 6953 7910 6958 7938
rect 6986 7910 7574 7938
rect 7602 7910 7607 7938
rect 10705 7910 10710 7938
rect 10738 7910 10990 7938
rect 11018 7910 11023 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 0 7770 400 7784
rect 20600 7770 21000 7784
rect 0 7742 1022 7770
rect 1050 7742 1055 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 0 7728 400 7742
rect 20600 7728 21000 7742
rect 8801 7686 8806 7714
rect 8834 7686 13230 7714
rect 13258 7686 13263 7714
rect 7737 7574 7742 7602
rect 7770 7574 8862 7602
rect 8890 7574 8895 7602
rect 9921 7574 9926 7602
rect 9954 7574 10822 7602
rect 10850 7574 10855 7602
rect 9025 7462 9030 7490
rect 9058 7462 9198 7490
rect 9226 7462 9231 7490
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 11433 7406 11438 7434
rect 11466 7406 11718 7434
rect 11746 7406 11751 7434
rect 9641 7350 9646 7378
rect 9674 7350 9982 7378
rect 10010 7350 12614 7378
rect 12642 7350 13174 7378
rect 13202 7350 13207 7378
rect 9809 7294 9814 7322
rect 9842 7294 10430 7322
rect 10458 7294 10463 7322
rect 11041 7294 11046 7322
rect 11074 7294 11382 7322
rect 11410 7294 11415 7322
rect 9753 7238 9758 7266
rect 9786 7238 11102 7266
rect 11130 7238 11270 7266
rect 11298 7238 11303 7266
rect 11937 7238 11942 7266
rect 11970 7238 12670 7266
rect 12698 7238 12703 7266
rect 9249 7182 9254 7210
rect 9282 7182 10542 7210
rect 10570 7182 11718 7210
rect 11746 7182 11751 7210
rect 7569 7126 7574 7154
rect 7602 7126 8750 7154
rect 8778 7126 10374 7154
rect 10402 7126 10407 7154
rect 11433 7126 11438 7154
rect 11466 7126 11606 7154
rect 11634 7126 12390 7154
rect 12418 7126 12838 7154
rect 12866 7126 13118 7154
rect 13146 7126 13151 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 10873 6846 10878 6874
rect 10906 6846 11438 6874
rect 11466 6846 11471 6874
rect 9809 6790 9814 6818
rect 9842 6790 10150 6818
rect 10178 6790 10183 6818
rect 11041 6790 11046 6818
rect 11074 6790 12278 6818
rect 12306 6790 12311 6818
rect 9305 6734 9310 6762
rect 9338 6734 10598 6762
rect 10626 6734 10631 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8745 2030 8750 2058
rect 8778 2030 9254 2058
rect 9282 2030 9287 2058
rect 10089 2030 10094 2058
rect 10122 2030 10710 2058
rect 10738 2030 10743 2058
rect 12441 2030 12446 2058
rect 12474 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 11769 1806 11774 1834
rect 11802 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6888 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9856 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10976 0 1 10976
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _115_
timestamp 1698175906
transform -1 0 11760 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform -1 0 8624 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9688 0 -1 10192
box -43 -43 1107 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _118_
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _119_
timestamp 1698175906
transform -1 0 11200 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9744 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _121_
timestamp 1698175906
transform 1 0 7336 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10304 0 -1 10192
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10864 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 9520 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 7336 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _127_
timestamp 1698175906
transform -1 0 12208 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7952 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 7448 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7168 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _131_
timestamp 1698175906
transform -1 0 6384 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _132_
timestamp 1698175906
transform 1 0 7504 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform 1 0 8176 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform 1 0 13664 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform -1 0 10976 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _136_
timestamp 1698175906
transform -1 0 10304 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _137_
timestamp 1698175906
transform 1 0 8120 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8680 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform 1 0 12880 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _140_
timestamp 1698175906
transform -1 0 9072 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform -1 0 9184 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _142_
timestamp 1698175906
transform 1 0 13216 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _143_
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8400 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _145_
timestamp 1698175906
transform -1 0 9128 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8512 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7952 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 11760
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8904 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _150_
timestamp 1698175906
transform -1 0 8568 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _151_
timestamp 1698175906
transform -1 0 7168 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _152_
timestamp 1698175906
transform -1 0 6440 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform -1 0 11984 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698175906
transform 1 0 10024 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _155_
timestamp 1698175906
transform 1 0 9856 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _156_
timestamp 1698175906
transform -1 0 11368 0 1 9408
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _157_
timestamp 1698175906
transform 1 0 10640 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _158_
timestamp 1698175906
transform 1 0 13048 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13048 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 10136 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _161_
timestamp 1698175906
transform -1 0 11312 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _163_
timestamp 1698175906
transform 1 0 12824 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _164_
timestamp 1698175906
transform 1 0 8904 0 -1 11760
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _165_
timestamp 1698175906
transform -1 0 14000 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _166_
timestamp 1698175906
transform 1 0 14000 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _167_
timestamp 1698175906
transform -1 0 8848 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform -1 0 11592 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _169_
timestamp 1698175906
transform -1 0 11144 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _170_
timestamp 1698175906
transform 1 0 8064 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform -1 0 8288 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _172_
timestamp 1698175906
transform 1 0 7224 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _173_
timestamp 1698175906
transform 1 0 8960 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform 1 0 9800 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _175_
timestamp 1698175906
transform -1 0 10472 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _176_
timestamp 1698175906
transform 1 0 9968 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _177_
timestamp 1698175906
transform -1 0 9912 0 1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _178_
timestamp 1698175906
transform -1 0 12768 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11144 0 -1 13328
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _180_
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _181_
timestamp 1698175906
transform 1 0 8624 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _182_
timestamp 1698175906
transform 1 0 12880 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform 1 0 10808 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _184_
timestamp 1698175906
transform 1 0 11368 0 1 9408
box -43 -43 1107 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _185_
timestamp 1698175906
transform -1 0 11872 0 -1 9408
box -43 -43 2115 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _186_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11592 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _187_
timestamp 1698175906
transform 1 0 12208 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _188_
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform 1 0 13160 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _190_
timestamp 1698175906
transform -1 0 12432 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_
timestamp 1698175906
transform -1 0 11368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _193_
timestamp 1698175906
transform -1 0 11032 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _194_
timestamp 1698175906
transform -1 0 11760 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _195_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9352 0 -1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _196_
timestamp 1698175906
transform 1 0 9464 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698175906
transform -1 0 9464 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _198_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10360 0 1 9408
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _199_
timestamp 1698175906
transform 1 0 13496 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1698175906
transform -1 0 13440 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _201_
timestamp 1698175906
transform 1 0 9016 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform 1 0 7168 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _203_
timestamp 1698175906
transform 1 0 8400 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _204_
timestamp 1698175906
transform 1 0 7448 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _205_
timestamp 1698175906
transform 1 0 8904 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _206_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9352 0 -1 7840
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _207_
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _208_
timestamp 1698175906
transform -1 0 12040 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform -1 0 12824 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _210_
timestamp 1698175906
transform -1 0 11592 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _211_
timestamp 1698175906
transform -1 0 12376 0 -1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _212_
timestamp 1698175906
transform -1 0 9520 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _213_
timestamp 1698175906
transform 1 0 7224 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _214_
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _215_
timestamp 1698175906
transform 1 0 7280 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _216_
timestamp 1698175906
transform 1 0 7616 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _217_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10080 0 1 11760
box -43 -43 995 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _218_
timestamp 1698175906
transform 1 0 9912 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _219_
timestamp 1698175906
transform 1 0 10248 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11480 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform -1 0 6552 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 12936 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 10920 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 6384 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 5656 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 5432 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 12768 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 13328 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 7000 0 1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 8960 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 11368 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 7000 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 10752 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 12768 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform -1 0 7448 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 7280 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 11312 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 11592 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform -1 0 7280 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform -1 0 7392 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 8848 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _247_
timestamp 1698175906
transform 1 0 13832 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _248_
timestamp 1698175906
transform 1 0 14560 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _249_
timestamp 1698175906
transform 1 0 14896 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 6776 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 12824 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 7896 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 7392 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 7168 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 14616 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 13440 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 9072 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 8848 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 13104 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 9184 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 12376 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 14504 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 12320 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 10360 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 14504 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 7560 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 8904 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform -1 0 13160 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 14056 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 8232 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 7504 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform -1 0 8848 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 8792 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9520 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11088 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11592 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 12040 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 8456 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_143
timestamp 1698175906
transform 1 0 8680 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_185
timestamp 1698175906
transform 1 0 11032 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_189
timestamp 1698175906
transform 1 0 11256 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_219
timestamp 1698175906
transform 1 0 12936 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_223 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13160 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698175906
transform 1 0 14056 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698175906
transform 1 0 14280 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_88
timestamp 1698175906
transform 1 0 5600 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_121
timestamp 1698175906
transform 1 0 7448 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_125
timestamp 1698175906
transform 1 0 7672 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_133
timestamp 1698175906
transform 1 0 8120 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_137
timestamp 1698175906
transform 1 0 8344 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698175906
transform 1 0 8456 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_179
timestamp 1698175906
transform 1 0 10696 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_218
timestamp 1698175906
transform 1 0 12880 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_250
timestamp 1698175906
transform 1 0 14672 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_266
timestamp 1698175906
transform 1 0 15568 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698175906
transform 1 0 16016 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698175906
transform 1 0 16240 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_117
timestamp 1698175906
transform 1 0 7224 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_203
timestamp 1698175906
transform 1 0 12040 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_207
timestamp 1698175906
transform 1 0 12264 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_211
timestamp 1698175906
transform 1 0 12488 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_219
timestamp 1698175906
transform 1 0 12936 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_221
timestamp 1698175906
transform 1 0 13048 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_228
timestamp 1698175906
transform 1 0 13440 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_88
timestamp 1698175906
transform 1 0 5600 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_90
timestamp 1698175906
transform 1 0 5712 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_120
timestamp 1698175906
transform 1 0 7392 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_124
timestamp 1698175906
transform 1 0 7616 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_155
timestamp 1698175906
transform 1 0 9352 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_163
timestamp 1698175906
transform 1 0 9800 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_193
timestamp 1698175906
transform 1 0 11480 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_197
timestamp 1698175906
transform 1 0 11704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_205
timestamp 1698175906
transform 1 0 12152 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_245
timestamp 1698175906
transform 1 0 14392 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_249
timestamp 1698175906
transform 1 0 14616 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_265
timestamp 1698175906
transform 1 0 15512 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_273
timestamp 1698175906
transform 1 0 15960 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 2464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_115
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_129
timestamp 1698175906
transform 1 0 7896 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_145
timestamp 1698175906
transform 1 0 8792 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_149
timestamp 1698175906
transform 1 0 9016 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_165
timestamp 1698175906
transform 1 0 9912 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 10360 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 11032 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_189
timestamp 1698175906
transform 1 0 11256 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_198
timestamp 1698175906
transform 1 0 11760 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_214
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_222
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_226
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_228
timestamp 1698175906
transform 1 0 13440 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_235
timestamp 1698175906
transform 1 0 13832 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 14280 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_123
timestamp 1698175906
transform 1 0 7560 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_133
timestamp 1698175906
transform 1 0 8120 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 8344 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698175906
transform 1 0 8848 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_148
timestamp 1698175906
transform 1 0 8960 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_155
timestamp 1698175906
transform 1 0 9352 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_171
timestamp 1698175906
transform 1 0 10248 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_175
timestamp 1698175906
transform 1 0 10472 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_182
timestamp 1698175906
transform 1 0 10864 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_198
timestamp 1698175906
transform 1 0 11760 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 12208 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_216
timestamp 1698175906
transform 1 0 12768 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_248
timestamp 1698175906
transform 1 0 14560 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698175906
transform 1 0 7112 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_122
timestamp 1698175906
transform 1 0 7504 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_132
timestamp 1698175906
transform 1 0 8064 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_136
timestamp 1698175906
transform 1 0 8288 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 10304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_237
timestamp 1698175906
transform 1 0 13944 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 14168 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_118
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_122
timestamp 1698175906
transform 1 0 7504 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698175906
transform 1 0 8400 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_158
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_162
timestamp 1698175906
transform 1 0 9744 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_217
timestamp 1698175906
transform 1 0 12824 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_223
timestamp 1698175906
transform 1 0 13160 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_225
timestamp 1698175906
transform 1 0 13272 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_255
timestamp 1698175906
transform 1 0 14952 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_271
timestamp 1698175906
transform 1 0 15848 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_131
timestamp 1698175906
transform 1 0 8008 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_147
timestamp 1698175906
transform 1 0 8904 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_226
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_260
timestamp 1698175906
transform 1 0 15232 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_292
timestamp 1698175906
transform 1 0 17024 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 17920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 18144 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 18256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_112
timestamp 1698175906
transform 1 0 6944 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_127
timestamp 1698175906
transform 1 0 7784 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 8288 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_161
timestamp 1698175906
transform 1 0 9688 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_163
timestamp 1698175906
transform 1 0 9800 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 16128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_236
timestamp 1698175906
transform 1 0 13888 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_84
timestamp 1698175906
transform 1 0 5376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_114
timestamp 1698175906
transform 1 0 7056 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_118
timestamp 1698175906
transform 1 0 7280 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_155
timestamp 1698175906
transform 1 0 9352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_157
timestamp 1698175906
transform 1 0 9464 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 12320 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_225
timestamp 1698175906
transform 1 0 13272 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_257
timestamp 1698175906
transform 1 0 15064 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698175906
transform 1 0 15960 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 16184 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_69
timestamp 1698175906
transform 1 0 4536 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_85
timestamp 1698175906
transform 1 0 5432 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_93
timestamp 1698175906
transform 1 0 5880 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698175906
transform 1 0 6440 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_116
timestamp 1698175906
transform 1 0 7168 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_132
timestamp 1698175906
transform 1 0 8064 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_141
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_251
timestamp 1698175906
transform 1 0 14728 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_96
timestamp 1698175906
transform 1 0 6048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_102
timestamp 1698175906
transform 1 0 6384 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_121
timestamp 1698175906
transform 1 0 7448 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_129
timestamp 1698175906
transform 1 0 7896 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_133
timestamp 1698175906
transform 1 0 8120 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698175906
transform 1 0 8736 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_195
timestamp 1698175906
transform 1 0 11592 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_245
timestamp 1698175906
transform 1 0 14392 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_249
timestamp 1698175906
transform 1 0 14616 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_265
timestamp 1698175906
transform 1 0 15512 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 15960 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_69
timestamp 1698175906
transform 1 0 4536 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_73
timestamp 1698175906
transform 1 0 4760 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_75
timestamp 1698175906
transform 1 0 4872 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_111
timestamp 1698175906
transform 1 0 6888 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_119
timestamp 1698175906
transform 1 0 7336 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_123
timestamp 1698175906
transform 1 0 7560 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_168
timestamp 1698175906
transform 1 0 10080 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_181
timestamp 1698175906
transform 1 0 10808 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_188
timestamp 1698175906
transform 1 0 11200 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_204
timestamp 1698175906
transform 1 0 12096 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_212
timestamp 1698175906
transform 1 0 12544 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_216
timestamp 1698175906
transform 1 0 12768 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_228
timestamp 1698175906
transform 1 0 13440 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_232
timestamp 1698175906
transform 1 0 13664 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_234
timestamp 1698175906
transform 1 0 13776 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_96
timestamp 1698175906
transform 1 0 6048 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_100
timestamp 1698175906
transform 1 0 6272 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_131
timestamp 1698175906
transform 1 0 8008 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_133
timestamp 1698175906
transform 1 0 8120 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_150
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_162
timestamp 1698175906
transform 1 0 9744 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_166
timestamp 1698175906
transform 1 0 9968 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_173
timestamp 1698175906
transform 1 0 10360 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_189
timestamp 1698175906
transform 1 0 11256 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 12208 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 16128 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_127
timestamp 1698175906
transform 1 0 7784 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_142
timestamp 1698175906
transform 1 0 8624 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_144
timestamp 1698175906
transform 1 0 8736 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_151
timestamp 1698175906
transform 1 0 9128 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_159
timestamp 1698175906
transform 1 0 9576 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698175906
transform 1 0 10080 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 10304 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_182
timestamp 1698175906
transform 1 0 10864 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_212
timestamp 1698175906
transform 1 0 12544 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_216
timestamp 1698175906
transform 1 0 12768 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_232
timestamp 1698175906
transform 1 0 13664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698175906
transform 1 0 14112 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_151
timestamp 1698175906
transform 1 0 9128 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_167
timestamp 1698175906
transform 1 0 10024 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_175
timestamp 1698175906
transform 1 0 10472 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_179
timestamp 1698175906
transform 1 0 10696 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_199
timestamp 1698175906
transform 1 0 11816 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 12264 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_216
timestamp 1698175906
transform 1 0 12768 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_150
timestamp 1698175906
transform 1 0 9072 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_154
timestamp 1698175906
transform 1 0 9296 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_165
timestamp 1698175906
transform 1 0 9912 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 10416 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698175906
transform 1 0 11032 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_189
timestamp 1698175906
transform 1 0 11256 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_220
timestamp 1698175906
transform 1 0 12992 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_224
timestamp 1698175906
transform 1 0 13216 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_240
timestamp 1698175906
transform 1 0 14112 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 7392 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_128
timestamp 1698175906
transform 1 0 7840 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_146
timestamp 1698175906
transform 1 0 8848 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_185
timestamp 1698175906
transform 1 0 11032 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_191
timestamp 1698175906
transform 1 0 11368 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 12264 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_111
timestamp 1698175906
transform 1 0 6888 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_142
timestamp 1698175906
transform 1 0 8624 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_148
timestamp 1698175906
transform 1 0 8960 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_152
timestamp 1698175906
transform 1 0 9184 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_168
timestamp 1698175906
transform 1 0 10080 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 10304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 10416 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_206
timestamp 1698175906
transform 1 0 12208 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_210
timestamp 1698175906
transform 1 0 12432 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 14336 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_333
timestamp 1698175906
transform 1 0 19320 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_341
timestamp 1698175906
transform 1 0 19768 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_172
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_204
timestamp 1698175906
transform 1 0 12096 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698175906
transform 1 0 12320 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 14280 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 16072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 10416 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 11928 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 12040 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita20_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10304 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita20_26
timestamp 1698175906
transform 1 0 19992 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 10136 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 2240 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 8680 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 10192 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 12824 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 10472 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 14112 400 14168 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 17136 21000 17192 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 7728 400 7784 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 11424 20600 11480 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 11732 13468 11732 13468 0 _000_
rlabel metal3 8120 13468 8120 13468 0 _001_
rlabel metal2 11228 7056 11228 7056 0 _002_
rlabel metal3 12768 11508 12768 11508 0 _003_
rlabel metal2 10892 14168 10892 14168 0 _004_
rlabel metal2 9100 7112 9100 7112 0 _005_
rlabel metal2 13244 7448 13244 7448 0 _006_
rlabel metal2 6972 7420 6972 7420 0 _007_
rlabel metal3 8316 7588 8316 7588 0 _008_
rlabel metal2 11732 6524 11732 6524 0 _009_
rlabel metal2 12096 8876 12096 8876 0 _010_
rlabel metal2 6804 8568 6804 8568 0 _011_
rlabel metal2 6916 8036 6916 8036 0 _012_
rlabel metal2 9324 6636 9324 6636 0 _013_
rlabel metal2 11004 7812 11004 7812 0 _014_
rlabel metal2 6244 11788 6244 11788 0 _015_
rlabel metal2 13384 8484 13384 8484 0 _016_
rlabel metal3 11900 11116 11900 11116 0 _017_
rlabel metal2 8260 12152 8260 12152 0 _018_
rlabel metal2 6132 9352 6132 9352 0 _019_
rlabel metal2 5908 10948 5908 10948 0 _020_
rlabel metal2 13216 11228 13216 11228 0 _021_
rlabel metal2 13804 9296 13804 9296 0 _022_
rlabel metal2 8204 14140 8204 14140 0 _023_
rlabel metal2 9548 13720 9548 13720 0 _024_
rlabel metal2 12992 11844 12992 11844 0 _025_
rlabel metal2 11228 11732 11228 11732 0 _026_
rlabel metal2 11172 11928 11172 11928 0 _027_
rlabel metal2 12124 11732 12124 11732 0 _028_
rlabel metal2 13636 9324 13636 9324 0 _029_
rlabel metal2 13972 9660 13972 9660 0 _030_
rlabel metal3 8484 13916 8484 13916 0 _031_
rlabel metal2 11564 12460 11564 12460 0 _032_
rlabel metal2 10920 13916 10920 13916 0 _033_
rlabel metal3 9100 13524 9100 13524 0 _034_
rlabel metal3 10444 9660 10444 9660 0 _035_
rlabel metal2 9604 12348 9604 12348 0 _036_
rlabel metal2 9940 12936 9940 12936 0 _037_
rlabel metal2 10220 11144 10220 11144 0 _038_
rlabel metal2 9968 13524 9968 13524 0 _039_
rlabel metal3 12152 13132 12152 13132 0 _040_
rlabel metal2 8932 13482 8932 13482 0 _041_
rlabel metal3 11844 8428 11844 8428 0 _042_
rlabel metal3 11228 7308 11228 7308 0 _043_
rlabel metal2 11508 9492 11508 9492 0 _044_
rlabel via2 11452 7420 11452 7420 0 _045_
rlabel metal2 12376 11060 12376 11060 0 _046_
rlabel metal2 12460 9492 12460 9492 0 _047_
rlabel metal2 12404 11704 12404 11704 0 _048_
rlabel metal3 11032 13916 11032 13916 0 _049_
rlabel metal2 10724 13412 10724 13412 0 _050_
rlabel metal2 11564 7924 11564 7924 0 _051_
rlabel metal2 9212 11424 9212 11424 0 _052_
rlabel metal2 9492 7308 9492 7308 0 _053_
rlabel metal3 9660 9464 9660 9464 0 _054_
rlabel metal2 13636 7756 13636 7756 0 _055_
rlabel metal2 9268 8428 9268 8428 0 _056_
rlabel metal2 7476 7980 7476 7980 0 _057_
rlabel metal2 8960 7644 8960 7644 0 _058_
rlabel metal2 9240 7644 9240 7644 0 _059_
rlabel metal2 12684 7112 12684 7112 0 _060_
rlabel metal2 12572 9184 12572 9184 0 _061_
rlabel metal2 11452 9072 11452 9072 0 _062_
rlabel metal2 7980 8848 7980 8848 0 _063_
rlabel metal3 7616 8708 7616 8708 0 _064_
rlabel metal3 7672 8428 7672 8428 0 _065_
rlabel metal2 9912 8708 9912 8708 0 _066_
rlabel metal2 10332 7084 10332 7084 0 _067_
rlabel metal2 11340 11060 11340 11060 0 _068_
rlabel metal2 7140 10248 7140 10248 0 _069_
rlabel metal2 11144 9996 11144 9996 0 _070_
rlabel metal2 10220 11564 10220 11564 0 _071_
rlabel metal3 10948 8540 10948 8540 0 _072_
rlabel metal2 8316 11872 8316 11872 0 _073_
rlabel metal2 8792 12236 8792 12236 0 _074_
rlabel metal2 10668 9100 10668 9100 0 _075_
rlabel metal2 10780 8820 10780 8820 0 _076_
rlabel metal2 12292 9800 12292 9800 0 _077_
rlabel metal2 10892 10220 10892 10220 0 _078_
rlabel metal2 7252 9968 7252 9968 0 _079_
rlabel metal2 10500 9688 10500 9688 0 _080_
rlabel metal2 10780 8456 10780 8456 0 _081_
rlabel metal2 7308 11648 7308 11648 0 _082_
rlabel metal2 6916 10850 6916 10850 0 _083_
rlabel metal2 8596 11872 8596 11872 0 _084_
rlabel metal2 8708 11200 8708 11200 0 _085_
rlabel metal3 7028 11676 7028 11676 0 _086_
rlabel metal3 6664 11564 6664 11564 0 _087_
rlabel metal2 8848 11172 8848 11172 0 _088_
rlabel metal2 13916 10822 13916 10822 0 _089_
rlabel metal3 13692 8764 13692 8764 0 _090_
rlabel metal2 12124 9856 12124 9856 0 _091_
rlabel metal2 9044 11368 9044 11368 0 _092_
rlabel metal2 10780 9856 10780 9856 0 _093_
rlabel metal2 13244 8260 13244 8260 0 _094_
rlabel metal2 8680 9212 8680 9212 0 _095_
rlabel metal2 13524 8848 13524 8848 0 _096_
rlabel metal3 9800 12684 9800 12684 0 _097_
rlabel metal2 8820 9660 8820 9660 0 _098_
rlabel metal2 8344 12348 8344 12348 0 _099_
rlabel metal3 8316 11956 8316 11956 0 _100_
rlabel metal2 8484 13678 8484 13678 0 _101_
rlabel metal3 7700 11172 7700 11172 0 _102_
rlabel metal3 6580 11116 6580 11116 0 _103_
rlabel metal2 12628 9576 12628 9576 0 _104_
rlabel metal2 10192 13468 10192 13468 0 _105_
rlabel metal2 11172 9548 11172 9548 0 _106_
rlabel metal3 11900 9604 11900 9604 0 _107_
rlabel metal2 10836 10500 10836 10500 0 _108_
rlabel metal2 13188 11004 13188 11004 0 _109_
rlabel metal3 1239 14140 1239 14140 0 clk
rlabel metal2 11172 10556 11172 10556 0 clknet_0_clk
rlabel metal3 6384 10780 6384 10780 0 clknet_1_0__leaf_clk
rlabel metal2 11452 13888 11452 13888 0 clknet_1_1__leaf_clk
rlabel metal3 12292 12460 12292 12460 0 dut20.count\[0\]
rlabel metal2 10164 12180 10164 12180 0 dut20.count\[1\]
rlabel metal2 7308 9772 7308 9772 0 dut20.count\[2\]
rlabel metal2 6972 10556 6972 10556 0 dut20.count\[3\]
rlabel metal3 15960 9184 15960 9184 0 net1
rlabel metal2 8988 4676 8988 4676 0 net10
rlabel metal2 12852 4340 12852 4340 0 net11
rlabel metal2 12292 4284 12292 4284 0 net12
rlabel metal2 8540 13692 8540 13692 0 net13
rlabel metal3 9996 6804 9996 6804 0 net14
rlabel metal2 14308 7812 14308 7812 0 net15
rlabel metal2 12796 13580 12796 13580 0 net16
rlabel metal2 10388 13692 10388 13692 0 net17
rlabel metal2 8764 14168 8764 14168 0 net18
rlabel metal2 18788 9744 18788 9744 0 net19
rlabel metal2 5740 8596 5740 8596 0 net2
rlabel metal2 14308 11032 14308 11032 0 net20
rlabel metal2 14476 8596 14476 8596 0 net21
rlabel metal3 3178 11956 3178 11956 0 net22
rlabel metal3 11704 13972 11704 13972 0 net23
rlabel metal3 10948 7980 10948 7980 0 net24
rlabel metal2 10164 19012 10164 19012 0 net25
rlabel metal2 20132 17248 20132 17248 0 net26
rlabel metal2 5852 8008 5852 8008 0 net3
rlabel metal2 10388 4340 10388 4340 0 net4
rlabel metal2 18844 11704 18844 11704 0 net5
rlabel metal2 14812 9576 14812 9576 0 net6
rlabel metal2 14308 11732 14308 11732 0 net7
rlabel metal2 15036 9576 15036 9576 0 net8
rlabel metal2 5908 7420 5908 7420 0 net9
rlabel metal3 20321 9100 20321 9100 0 segm[10]
rlabel metal3 679 8764 679 8764 0 segm[11]
rlabel metal3 679 8092 679 8092 0 segm[12]
rlabel metal3 10416 2044 10416 2044 0 segm[13]
rlabel metal3 20321 11452 20321 11452 0 segm[1]
rlabel metal2 20020 10276 20020 10276 0 segm[2]
rlabel metal2 20020 11900 20020 11900 0 segm[4]
rlabel metal2 20020 9548 20020 9548 0 segm[5]
rlabel metal3 707 7756 707 7756 0 segm[6]
rlabel metal3 9016 2044 9016 2044 0 segm[7]
rlabel metal3 12796 2044 12796 2044 0 segm[8]
rlabel metal3 12292 1820 12292 1820 0 segm[9]
rlabel metal2 8428 19677 8428 19677 0 sel[0]
rlabel metal2 9772 1015 9772 1015 0 sel[10]
rlabel metal2 20020 7924 20020 7924 0 sel[11]
rlabel metal2 12796 19957 12796 19957 0 sel[1]
rlabel metal2 10444 19873 10444 19873 0 sel[2]
rlabel metal2 8764 19873 8764 19873 0 sel[3]
rlabel metal2 20020 9828 20020 9828 0 sel[4]
rlabel metal2 20020 11172 20020 11172 0 sel[5]
rlabel metal2 20020 8820 20020 8820 0 sel[6]
rlabel metal3 679 11788 679 11788 0 sel[7]
rlabel metal2 11452 19873 11452 19873 0 sel[8]
rlabel metal2 11116 1015 11116 1015 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
