magic
tech gf180mcuD
magscale 1 5
timestamp 1699644056
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9591 19137 9617 19143
rect 9591 19105 9617 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9865 18999 9871 19025
rect 9897 18999 9903 19025
rect 10705 18999 10711 19025
rect 10737 18999 10743 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 13735 18969 13761 18975
rect 13735 18937 13761 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9367 18745 9393 18751
rect 9367 18713 9393 18719
rect 11047 18745 11073 18751
rect 11047 18713 11073 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 8857 18607 8863 18633
rect 8889 18607 8895 18633
rect 10649 18607 10655 18633
rect 10681 18607 10687 18633
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 13399 18353 13425 18359
rect 13399 18321 13425 18327
rect 12889 18215 12895 18241
rect 12921 18215 12927 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 9927 14433 9953 14439
rect 9927 14401 9953 14407
rect 11663 14433 11689 14439
rect 11663 14401 11689 14407
rect 12217 14295 12223 14321
rect 12249 14295 12255 14321
rect 9983 14265 10009 14271
rect 9983 14233 10009 14239
rect 10207 14265 10233 14271
rect 10207 14233 10233 14239
rect 10263 14265 10289 14271
rect 10263 14233 10289 14239
rect 11607 14265 11633 14271
rect 12329 14239 12335 14265
rect 12361 14239 12367 14265
rect 11607 14233 11633 14239
rect 9927 14209 9953 14215
rect 9927 14177 9953 14183
rect 10095 14209 10121 14215
rect 10095 14177 10121 14183
rect 11663 14209 11689 14215
rect 11663 14177 11689 14183
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 12671 14041 12697 14047
rect 12671 14009 12697 14015
rect 9585 13959 9591 13985
rect 9617 13959 9623 13985
rect 11265 13959 11271 13985
rect 11297 13959 11303 13985
rect 12615 13929 12641 13935
rect 9249 13903 9255 13929
rect 9281 13903 9287 13929
rect 10873 13903 10879 13929
rect 10905 13903 10911 13929
rect 12615 13897 12641 13903
rect 13007 13929 13033 13935
rect 13007 13897 13033 13903
rect 10649 13847 10655 13873
rect 10681 13847 10687 13873
rect 12329 13847 12335 13873
rect 12361 13847 12367 13873
rect 12671 13817 12697 13823
rect 12671 13785 12697 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10767 13593 10793 13599
rect 13119 13593 13145 13599
rect 9977 13567 9983 13593
rect 10009 13567 10015 13593
rect 12889 13567 12895 13593
rect 12921 13567 12927 13593
rect 10767 13561 10793 13567
rect 13119 13561 13145 13567
rect 8359 13537 8385 13543
rect 10151 13537 10177 13543
rect 8521 13511 8527 13537
rect 8553 13511 8559 13537
rect 11433 13511 11439 13537
rect 11465 13511 11471 13537
rect 8359 13505 8385 13511
rect 10151 13505 10177 13511
rect 10263 13481 10289 13487
rect 8913 13455 8919 13481
rect 8945 13455 8951 13481
rect 10263 13449 10289 13455
rect 10319 13481 10345 13487
rect 11825 13455 11831 13481
rect 11857 13455 11863 13481
rect 10319 13449 10345 13455
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 9143 13257 9169 13263
rect 11551 13257 11577 13263
rect 10313 13231 10319 13257
rect 10345 13231 10351 13257
rect 9143 13225 9169 13231
rect 11551 13225 11577 13231
rect 11663 13257 11689 13263
rect 11663 13225 11689 13231
rect 11831 13257 11857 13263
rect 11831 13225 11857 13231
rect 8751 13201 8777 13207
rect 8751 13169 8777 13175
rect 9255 13201 9281 13207
rect 9255 13169 9281 13175
rect 9311 13201 9337 13207
rect 9311 13169 9337 13175
rect 11719 13201 11745 13207
rect 11719 13169 11745 13175
rect 11943 13201 11969 13207
rect 11943 13169 11969 13175
rect 11999 13201 12025 13207
rect 11999 13169 12025 13175
rect 10151 13145 10177 13151
rect 7009 13119 7015 13145
rect 7041 13119 7047 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 10151 13113 10177 13119
rect 7345 13063 7351 13089
rect 7377 13063 7383 13089
rect 8409 13063 8415 13089
rect 8441 13063 8447 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 967 12809 993 12815
rect 8527 12809 8553 12815
rect 4993 12783 4999 12809
rect 5025 12783 5031 12809
rect 967 12777 993 12783
rect 8527 12777 8553 12783
rect 20007 12809 20033 12815
rect 20007 12777 20033 12783
rect 8639 12753 8665 12759
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 6449 12727 6455 12753
rect 6481 12727 6487 12753
rect 8639 12721 8665 12727
rect 12783 12753 12809 12759
rect 12783 12721 12809 12727
rect 12951 12753 12977 12759
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 12951 12721 12977 12727
rect 6791 12697 6817 12703
rect 6057 12671 6063 12697
rect 6089 12671 6095 12697
rect 6791 12665 6817 12671
rect 7967 12697 7993 12703
rect 7967 12665 7993 12671
rect 8135 12697 8161 12703
rect 8135 12665 8161 12671
rect 10655 12697 10681 12703
rect 10655 12665 10681 12671
rect 13007 12697 13033 12703
rect 13007 12665 13033 12671
rect 6735 12641 6761 12647
rect 6735 12609 6761 12615
rect 7015 12641 7041 12647
rect 10711 12641 10737 12647
rect 8801 12615 8807 12641
rect 8833 12615 8839 12641
rect 7015 12609 7041 12615
rect 10711 12609 10737 12615
rect 10823 12641 10849 12647
rect 10823 12609 10849 12615
rect 12615 12641 12641 12647
rect 12615 12609 12641 12615
rect 12727 12641 12753 12647
rect 12727 12609 12753 12615
rect 13119 12641 13145 12647
rect 13119 12609 13145 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 8695 12473 8721 12479
rect 8695 12441 8721 12447
rect 12223 12473 12249 12479
rect 12223 12441 12249 12447
rect 6561 12391 6567 12417
rect 6593 12391 6599 12417
rect 14401 12391 14407 12417
rect 14433 12391 14439 12417
rect 9031 12361 9057 12367
rect 12055 12361 12081 12367
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 6953 12335 6959 12361
rect 6985 12335 6991 12361
rect 11265 12335 11271 12361
rect 11297 12335 11303 12361
rect 9031 12329 9057 12335
rect 12055 12329 12081 12335
rect 12111 12361 12137 12367
rect 12111 12329 12137 12335
rect 12335 12361 12361 12367
rect 12665 12335 12671 12361
rect 12697 12335 12703 12361
rect 14289 12335 14295 12361
rect 14321 12335 14327 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 12335 12329 12361 12335
rect 7183 12305 7209 12311
rect 5497 12279 5503 12305
rect 5529 12279 5535 12305
rect 7183 12273 7209 12279
rect 9143 12305 9169 12311
rect 11495 12305 11521 12311
rect 9809 12279 9815 12305
rect 9841 12279 9847 12305
rect 10873 12279 10879 12305
rect 10905 12279 10911 12305
rect 9143 12273 9169 12279
rect 11495 12273 11521 12279
rect 12391 12305 12417 12311
rect 14631 12305 14657 12311
rect 13001 12279 13007 12305
rect 13033 12279 13039 12305
rect 14065 12279 14071 12305
rect 14097 12279 14103 12305
rect 12391 12273 12417 12279
rect 14631 12273 14657 12279
rect 967 12249 993 12255
rect 967 12217 993 12223
rect 8919 12249 8945 12255
rect 8919 12217 8945 12223
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 6399 12081 6425 12087
rect 6399 12049 6425 12055
rect 967 12025 993 12031
rect 6897 11999 6903 12025
rect 6929 11999 6935 12025
rect 7569 11999 7575 12025
rect 7601 11999 7607 12025
rect 10873 11999 10879 12025
rect 10905 11999 10911 12025
rect 13393 11999 13399 12025
rect 13425 11999 13431 12025
rect 967 11993 993 11999
rect 6455 11969 6481 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 6455 11937 6481 11943
rect 6959 11969 6985 11975
rect 9143 11969 9169 11975
rect 9025 11943 9031 11969
rect 9057 11943 9063 11969
rect 6959 11937 6985 11943
rect 9143 11937 9169 11943
rect 9311 11969 9337 11975
rect 13623 11969 13649 11975
rect 10649 11943 10655 11969
rect 10681 11943 10687 11969
rect 11657 11943 11663 11969
rect 11689 11943 11695 11969
rect 11993 11943 11999 11969
rect 12025 11943 12031 11969
rect 9311 11937 9337 11943
rect 13623 11937 13649 11943
rect 7183 11913 7209 11919
rect 9255 11913 9281 11919
rect 8633 11887 8639 11913
rect 8665 11887 8671 11913
rect 7183 11881 7209 11887
rect 9255 11881 9281 11887
rect 9479 11913 9505 11919
rect 9479 11881 9505 11887
rect 11551 11913 11577 11919
rect 12329 11887 12335 11913
rect 12361 11887 12367 11913
rect 11551 11881 11577 11887
rect 6903 11857 6929 11863
rect 6903 11825 6929 11831
rect 7071 11857 7097 11863
rect 7071 11825 7097 11831
rect 9703 11857 9729 11863
rect 9703 11825 9729 11831
rect 10767 11857 10793 11863
rect 10767 11825 10793 11831
rect 10879 11857 10905 11863
rect 10879 11825 10905 11831
rect 11775 11857 11801 11863
rect 11775 11825 11801 11831
rect 11831 11857 11857 11863
rect 11831 11825 11857 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 6959 11689 6985 11695
rect 6959 11657 6985 11663
rect 8807 11689 8833 11695
rect 8807 11657 8833 11663
rect 8863 11689 8889 11695
rect 8863 11657 8889 11663
rect 9367 11689 9393 11695
rect 9367 11657 9393 11663
rect 10375 11689 10401 11695
rect 11999 11689 12025 11695
rect 11713 11663 11719 11689
rect 11745 11663 11751 11689
rect 10375 11657 10401 11663
rect 11999 11657 12025 11663
rect 9255 11633 9281 11639
rect 9255 11601 9281 11607
rect 9927 11633 9953 11639
rect 9927 11601 9953 11607
rect 6847 11577 6873 11583
rect 6847 11545 6873 11551
rect 6903 11577 6929 11583
rect 6903 11545 6929 11551
rect 7015 11577 7041 11583
rect 7015 11545 7041 11551
rect 7071 11577 7097 11583
rect 7071 11545 7097 11551
rect 8751 11577 8777 11583
rect 8751 11545 8777 11551
rect 8919 11577 8945 11583
rect 9199 11577 9225 11583
rect 9025 11551 9031 11577
rect 9057 11551 9063 11577
rect 8919 11545 8945 11551
rect 9199 11545 9225 11551
rect 9871 11577 9897 11583
rect 9871 11545 9897 11551
rect 10039 11577 10065 11583
rect 11887 11577 11913 11583
rect 10481 11551 10487 11577
rect 10513 11551 10519 11577
rect 12105 11551 12111 11577
rect 12137 11551 12143 11577
rect 12217 11551 12223 11577
rect 12249 11551 12255 11577
rect 10039 11545 10065 11551
rect 11887 11545 11913 11551
rect 10319 11521 10345 11527
rect 10319 11489 10345 11495
rect 11439 11521 11465 11527
rect 11439 11489 11465 11495
rect 11551 11521 11577 11527
rect 12671 11521 12697 11527
rect 12273 11495 12279 11521
rect 12305 11495 12311 11521
rect 11551 11489 11577 11495
rect 12671 11489 12697 11495
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 12559 11297 12585 11303
rect 12559 11265 12585 11271
rect 967 11241 993 11247
rect 20007 11241 20033 11247
rect 14233 11215 14239 11241
rect 14265 11215 14271 11241
rect 967 11209 993 11215
rect 20007 11209 20033 11215
rect 6735 11185 6761 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 6735 11153 6761 11159
rect 6959 11185 6985 11191
rect 6959 11153 6985 11159
rect 7183 11185 7209 11191
rect 7183 11153 7209 11159
rect 7351 11185 7377 11191
rect 8247 11185 8273 11191
rect 7961 11159 7967 11185
rect 7993 11159 7999 11185
rect 7351 11153 7377 11159
rect 8247 11153 8273 11159
rect 8919 11185 8945 11191
rect 8919 11153 8945 11159
rect 9143 11185 9169 11191
rect 11047 11185 11073 11191
rect 9585 11159 9591 11185
rect 9617 11159 9623 11185
rect 9809 11159 9815 11185
rect 9841 11159 9847 11185
rect 10257 11159 10263 11185
rect 10289 11159 10295 11185
rect 9143 11153 9169 11159
rect 11047 11153 11073 11159
rect 12279 11185 12305 11191
rect 12279 11153 12305 11159
rect 12503 11185 12529 11191
rect 12777 11159 12783 11185
rect 12809 11159 12815 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 12503 11153 12529 11159
rect 6903 11129 6929 11135
rect 11215 11129 11241 11135
rect 9473 11103 9479 11129
rect 9505 11103 9511 11129
rect 10313 11103 10319 11129
rect 10345 11103 10351 11129
rect 6903 11097 6929 11103
rect 11215 11097 11241 11103
rect 12615 11129 12641 11135
rect 13169 11103 13175 11129
rect 13201 11103 13207 11129
rect 12615 11097 12641 11103
rect 6791 11073 6817 11079
rect 6791 11041 6817 11047
rect 7239 11073 7265 11079
rect 8303 11073 8329 11079
rect 8073 11047 8079 11073
rect 8105 11047 8111 11073
rect 7239 11041 7265 11047
rect 8303 11041 8329 11047
rect 8751 11073 8777 11079
rect 8751 11041 8777 11047
rect 8975 11073 9001 11079
rect 11159 11073 11185 11079
rect 9865 11047 9871 11073
rect 9897 11047 9903 11073
rect 8975 11041 9001 11047
rect 11159 11041 11185 11047
rect 12391 11073 12417 11079
rect 12391 11041 12417 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 12279 10905 12305 10911
rect 11881 10879 11887 10905
rect 11913 10879 11919 10905
rect 12279 10873 12305 10879
rect 12671 10905 12697 10911
rect 12671 10873 12697 10879
rect 13119 10905 13145 10911
rect 13119 10873 13145 10879
rect 13231 10905 13257 10911
rect 13231 10873 13257 10879
rect 8857 10823 8863 10849
rect 8889 10823 8895 10849
rect 8415 10793 8441 10799
rect 12223 10793 12249 10799
rect 6337 10767 6343 10793
rect 6369 10767 6375 10793
rect 8745 10767 8751 10793
rect 8777 10767 8783 10793
rect 9249 10767 9255 10793
rect 9281 10767 9287 10793
rect 11993 10767 11999 10793
rect 12025 10767 12031 10793
rect 8415 10761 8441 10767
rect 12223 10761 12249 10767
rect 12391 10793 12417 10799
rect 12391 10761 12417 10767
rect 12783 10793 12809 10799
rect 12783 10761 12809 10767
rect 12895 10793 12921 10799
rect 12895 10761 12921 10767
rect 13063 10793 13089 10799
rect 13063 10761 13089 10767
rect 7967 10737 7993 10743
rect 12839 10737 12865 10743
rect 6673 10711 6679 10737
rect 6705 10711 6711 10737
rect 7737 10711 7743 10737
rect 7769 10711 7775 10737
rect 8185 10711 8191 10737
rect 8217 10711 8223 10737
rect 10817 10711 10823 10737
rect 10849 10711 10855 10737
rect 7967 10705 7993 10711
rect 12839 10705 12865 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 6791 10457 6817 10463
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 6057 10431 6063 10457
rect 6089 10431 6095 10457
rect 7961 10431 7967 10457
rect 7993 10431 7999 10457
rect 10033 10431 10039 10457
rect 10065 10431 10071 10457
rect 6791 10425 6817 10431
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 9809 10375 9815 10401
rect 9841 10375 9847 10401
rect 10201 10375 10207 10401
rect 10233 10375 10239 10401
rect 10817 10375 10823 10401
rect 10849 10375 10855 10401
rect 12833 10319 12839 10345
rect 12865 10319 12871 10345
rect 9983 10289 10009 10295
rect 9983 10257 10009 10263
rect 10095 10289 10121 10295
rect 10095 10257 10121 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 6791 10065 6817 10071
rect 6791 10033 6817 10039
rect 6959 10065 6985 10071
rect 6959 10033 6985 10039
rect 7071 10065 7097 10071
rect 7071 10033 7097 10039
rect 7351 10065 7377 10071
rect 7351 10033 7377 10039
rect 8695 10065 8721 10071
rect 8695 10033 8721 10039
rect 10375 10065 10401 10071
rect 11103 10065 11129 10071
rect 10705 10039 10711 10065
rect 10737 10039 10743 10065
rect 10375 10033 10401 10039
rect 11103 10033 11129 10039
rect 11439 10065 11465 10071
rect 11439 10033 11465 10039
rect 11607 10065 11633 10071
rect 11769 10039 11775 10065
rect 11801 10039 11807 10065
rect 13841 10039 13847 10065
rect 13873 10039 13879 10065
rect 11607 10033 11633 10039
rect 6903 10009 6929 10015
rect 6903 9977 6929 9983
rect 7015 10009 7041 10015
rect 10543 10009 10569 10015
rect 11271 10009 11297 10015
rect 7793 9983 7799 10009
rect 7825 9983 7831 10009
rect 8857 9983 8863 10009
rect 8889 9983 8895 10009
rect 9081 9983 9087 10009
rect 9113 9983 9119 10009
rect 9249 9983 9255 10009
rect 9281 9983 9287 10009
rect 9977 9983 9983 10009
rect 10009 9983 10015 10009
rect 10257 9983 10263 10009
rect 10289 9983 10295 10009
rect 10873 9983 10879 10009
rect 10905 9983 10911 10009
rect 10985 9983 10991 10009
rect 11017 9983 11023 10009
rect 12329 9983 12335 10009
rect 12361 9983 12367 10009
rect 14177 9983 14183 10009
rect 14209 9983 14215 10009
rect 7015 9977 7041 9983
rect 10543 9977 10569 9983
rect 11271 9977 11297 9983
rect 6511 9953 6537 9959
rect 7463 9953 7489 9959
rect 8135 9953 8161 9959
rect 7289 9927 7295 9953
rect 7321 9927 7327 9953
rect 7905 9927 7911 9953
rect 7937 9927 7943 9953
rect 6511 9921 6537 9927
rect 7463 9921 7489 9927
rect 8135 9921 8161 9927
rect 8751 9953 8777 9959
rect 8751 9921 8777 9927
rect 9759 9953 9785 9959
rect 9759 9921 9785 9927
rect 10935 9953 10961 9959
rect 12777 9927 12783 9953
rect 12809 9927 12815 9953
rect 10935 9921 10961 9927
rect 12167 9897 12193 9903
rect 9081 9871 9087 9897
rect 9113 9871 9119 9897
rect 12167 9865 12193 9871
rect 12335 9897 12361 9903
rect 12335 9865 12361 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 11047 9729 11073 9735
rect 7009 9703 7015 9729
rect 7041 9703 7047 9729
rect 11047 9697 11073 9703
rect 11439 9729 11465 9735
rect 11439 9697 11465 9703
rect 7183 9673 7209 9679
rect 5329 9647 5335 9673
rect 5361 9647 5367 9673
rect 6393 9647 6399 9673
rect 6425 9647 6431 9673
rect 7183 9641 7209 9647
rect 8807 9673 8833 9679
rect 20007 9673 20033 9679
rect 11209 9647 11215 9673
rect 11241 9647 11247 9673
rect 12049 9647 12055 9673
rect 12081 9647 12087 9673
rect 13225 9647 13231 9673
rect 13257 9647 13263 9673
rect 14289 9647 14295 9673
rect 14321 9647 14327 9673
rect 8807 9641 8833 9647
rect 20007 9641 20033 9647
rect 6735 9617 6761 9623
rect 4993 9591 4999 9617
rect 5025 9591 5031 9617
rect 6735 9585 6761 9591
rect 6847 9617 6873 9623
rect 6847 9585 6873 9591
rect 8023 9617 8049 9623
rect 8023 9585 8049 9591
rect 8471 9617 8497 9623
rect 8471 9585 8497 9591
rect 8695 9617 8721 9623
rect 8695 9585 8721 9591
rect 8919 9617 8945 9623
rect 8919 9585 8945 9591
rect 9031 9617 9057 9623
rect 10767 9617 10793 9623
rect 9361 9591 9367 9617
rect 9393 9591 9399 9617
rect 9697 9591 9703 9617
rect 9729 9591 9735 9617
rect 9921 9591 9927 9617
rect 9953 9591 9959 9617
rect 10313 9591 10319 9617
rect 10345 9591 10351 9617
rect 9031 9585 9057 9591
rect 10767 9585 10793 9591
rect 11999 9617 12025 9623
rect 12329 9591 12335 9617
rect 12361 9591 12367 9617
rect 12833 9591 12839 9617
rect 12865 9591 12871 9617
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 11999 9585 12025 9591
rect 7239 9561 7265 9567
rect 7239 9529 7265 9535
rect 8079 9561 8105 9567
rect 11159 9561 11185 9567
rect 8297 9535 8303 9561
rect 8329 9535 8335 9561
rect 9641 9535 9647 9561
rect 9673 9535 9679 9561
rect 10369 9535 10375 9561
rect 10401 9535 10407 9561
rect 8079 9529 8105 9535
rect 11159 9529 11185 9535
rect 11383 9561 11409 9567
rect 11383 9529 11409 9535
rect 11775 9561 11801 9567
rect 12441 9535 12447 9561
rect 12473 9535 12479 9561
rect 11775 9529 11801 9535
rect 8191 9505 8217 9511
rect 10823 9505 10849 9511
rect 9249 9479 9255 9505
rect 9281 9479 9287 9505
rect 8191 9473 8217 9479
rect 10823 9473 10849 9479
rect 10935 9505 10961 9511
rect 10935 9473 10961 9479
rect 11439 9505 11465 9511
rect 11439 9473 11465 9479
rect 11887 9505 11913 9511
rect 11887 9473 11913 9479
rect 12055 9505 12081 9511
rect 12055 9473 12081 9479
rect 12671 9505 12697 9511
rect 12671 9473 12697 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 6287 9337 6313 9343
rect 8359 9337 8385 9343
rect 7177 9311 7183 9337
rect 7209 9311 7215 9337
rect 6287 9305 6313 9311
rect 8359 9305 8385 9311
rect 9143 9337 9169 9343
rect 9143 9305 9169 9311
rect 9591 9337 9617 9343
rect 9591 9305 9617 9311
rect 10431 9337 10457 9343
rect 10431 9305 10457 9311
rect 11327 9337 11353 9343
rect 11327 9305 11353 9311
rect 13007 9337 13033 9343
rect 13007 9305 13033 9311
rect 8415 9281 8441 9287
rect 8415 9249 8441 9255
rect 8695 9281 8721 9287
rect 8695 9249 8721 9255
rect 9535 9281 9561 9287
rect 9535 9249 9561 9255
rect 10151 9281 10177 9287
rect 10151 9249 10177 9255
rect 10823 9281 10849 9287
rect 10823 9249 10849 9255
rect 10879 9281 10905 9287
rect 12615 9281 12641 9287
rect 11489 9255 11495 9281
rect 11521 9255 11527 9281
rect 10879 9249 10905 9255
rect 12615 9249 12641 9255
rect 6455 9225 6481 9231
rect 7015 9225 7041 9231
rect 6561 9199 6567 9225
rect 6593 9199 6599 9225
rect 6455 9193 6481 9199
rect 7015 9193 7041 9199
rect 8807 9225 8833 9231
rect 8807 9193 8833 9199
rect 8975 9225 9001 9231
rect 8975 9193 9001 9199
rect 9087 9225 9113 9231
rect 9087 9193 9113 9199
rect 9367 9225 9393 9231
rect 9367 9193 9393 9199
rect 9759 9225 9785 9231
rect 10319 9225 10345 9231
rect 13231 9225 13257 9231
rect 9865 9199 9871 9225
rect 9897 9199 9903 9225
rect 12721 9199 12727 9225
rect 12753 9199 12759 9225
rect 12889 9199 12895 9225
rect 12921 9199 12927 9225
rect 13337 9199 13343 9225
rect 13369 9199 13375 9225
rect 18937 9199 18943 9225
rect 18969 9199 18975 9225
rect 9759 9193 9785 9199
rect 10319 9193 10345 9199
rect 13231 9193 13257 9199
rect 6007 9169 6033 9175
rect 6007 9137 6033 9143
rect 9311 9169 9337 9175
rect 12335 9169 12361 9175
rect 10481 9143 10487 9169
rect 10513 9143 10519 9169
rect 9311 9137 9337 9143
rect 12335 9137 12361 9143
rect 8359 9113 8385 9119
rect 6785 9087 6791 9113
rect 6817 9087 6823 9113
rect 8359 9081 8385 9087
rect 10879 9113 10905 9119
rect 13175 9113 13201 9119
rect 12889 9087 12895 9113
rect 12921 9087 12927 9113
rect 10879 9081 10905 9087
rect 13175 9081 13201 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 6063 8945 6089 8951
rect 6063 8913 6089 8919
rect 11047 8945 11073 8951
rect 11047 8913 11073 8919
rect 6119 8889 6145 8895
rect 20007 8889 20033 8895
rect 7009 8863 7015 8889
rect 7041 8863 7047 8889
rect 13225 8863 13231 8889
rect 13257 8863 13263 8889
rect 14289 8863 14295 8889
rect 14321 8863 14327 8889
rect 6119 8857 6145 8863
rect 20007 8857 20033 8863
rect 7295 8833 7321 8839
rect 6897 8807 6903 8833
rect 6929 8807 6935 8833
rect 7295 8801 7321 8807
rect 9927 8833 9953 8839
rect 9927 8801 9953 8807
rect 10991 8833 11017 8839
rect 12833 8807 12839 8833
rect 12865 8807 12871 8833
rect 14625 8807 14631 8833
rect 14657 8807 14663 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 10991 8801 11017 8807
rect 9983 8777 10009 8783
rect 6281 8751 6287 8777
rect 6313 8751 6319 8777
rect 9983 8745 10009 8751
rect 10767 8777 10793 8783
rect 10767 8745 10793 8751
rect 6455 8721 6481 8727
rect 6455 8689 6481 8695
rect 10095 8721 10121 8727
rect 10095 8689 10121 8695
rect 10599 8721 10625 8727
rect 10599 8689 10625 8695
rect 10711 8721 10737 8727
rect 10711 8689 10737 8695
rect 11047 8721 11073 8727
rect 11047 8689 11073 8695
rect 12671 8721 12697 8727
rect 14737 8695 14743 8721
rect 14769 8695 14775 8721
rect 12671 8689 12697 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 8303 8553 8329 8559
rect 8303 8521 8329 8527
rect 8975 8553 9001 8559
rect 8975 8521 9001 8527
rect 9759 8553 9785 8559
rect 9759 8521 9785 8527
rect 10151 8553 10177 8559
rect 10151 8521 10177 8527
rect 10207 8553 10233 8559
rect 10207 8521 10233 8527
rect 7463 8497 7489 8503
rect 8079 8497 8105 8503
rect 5833 8471 5839 8497
rect 5865 8471 5871 8497
rect 7625 8471 7631 8497
rect 7657 8471 7663 8497
rect 7463 8465 7489 8471
rect 8079 8465 8105 8471
rect 8919 8497 8945 8503
rect 11607 8497 11633 8503
rect 9585 8471 9591 8497
rect 9617 8471 9623 8497
rect 8919 8465 8945 8471
rect 11607 8465 11633 8471
rect 11887 8497 11913 8503
rect 11887 8465 11913 8471
rect 9087 8441 9113 8447
rect 5497 8415 5503 8441
rect 5529 8415 5535 8441
rect 8185 8415 8191 8441
rect 8217 8415 8223 8441
rect 8689 8415 8695 8441
rect 8721 8415 8727 8441
rect 9087 8409 9113 8415
rect 10319 8441 10345 8447
rect 11663 8441 11689 8447
rect 10425 8415 10431 8441
rect 10457 8415 10463 8441
rect 10319 8409 10345 8415
rect 11663 8409 11689 8415
rect 11775 8441 11801 8447
rect 11775 8409 11801 8415
rect 7127 8385 7153 8391
rect 10263 8385 10289 8391
rect 6897 8359 6903 8385
rect 6929 8359 6935 8385
rect 8913 8359 8919 8385
rect 8945 8359 8951 8385
rect 7127 8353 7153 8359
rect 10263 8353 10289 8359
rect 8135 8329 8161 8335
rect 8135 8297 8161 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 12727 8161 12753 8167
rect 12727 8129 12753 8135
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 8303 8049 8329 8055
rect 8303 8017 8329 8023
rect 8415 8049 8441 8055
rect 8415 8017 8441 8023
rect 8639 8049 8665 8055
rect 8639 8017 8665 8023
rect 10599 8049 10625 8055
rect 10599 8017 10625 8023
rect 12167 8049 12193 8055
rect 12391 8049 12417 8055
rect 12783 8049 12809 8055
rect 12273 8023 12279 8049
rect 12305 8023 12311 8049
rect 12441 8023 12447 8049
rect 12473 8023 12479 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 12167 8017 12193 8023
rect 12391 8017 12417 8023
rect 12783 8017 12809 8023
rect 10711 7993 10737 7999
rect 10711 7961 10737 7967
rect 10767 7993 10793 7999
rect 10767 7961 10793 7967
rect 8359 7937 8385 7943
rect 8359 7905 8385 7911
rect 10991 7937 11017 7943
rect 10991 7905 11017 7911
rect 12559 7937 12585 7943
rect 12559 7905 12585 7911
rect 12839 7937 12865 7943
rect 12839 7905 12865 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8863 7769 8889 7775
rect 8863 7737 8889 7743
rect 9031 7769 9057 7775
rect 9031 7737 9057 7743
rect 12167 7769 12193 7775
rect 12167 7737 12193 7743
rect 14295 7769 14321 7775
rect 14295 7737 14321 7743
rect 8919 7713 8945 7719
rect 11159 7713 11185 7719
rect 7345 7687 7351 7713
rect 7377 7687 7383 7713
rect 9753 7687 9759 7713
rect 9785 7687 9791 7713
rect 8919 7681 8945 7687
rect 11159 7681 11185 7687
rect 11271 7713 11297 7719
rect 11271 7681 11297 7687
rect 11887 7713 11913 7719
rect 11887 7681 11913 7687
rect 12279 7713 12305 7719
rect 12279 7681 12305 7687
rect 12335 7713 12361 7719
rect 13001 7687 13007 7713
rect 13033 7687 13039 7713
rect 12335 7681 12361 7687
rect 9199 7657 9225 7663
rect 10935 7657 10961 7663
rect 7009 7631 7015 7657
rect 7041 7631 7047 7657
rect 9417 7631 9423 7657
rect 9449 7631 9455 7657
rect 9199 7625 9225 7631
rect 10935 7625 10961 7631
rect 11663 7657 11689 7663
rect 11663 7625 11689 7631
rect 11999 7657 12025 7663
rect 12609 7631 12615 7657
rect 12641 7631 12647 7657
rect 11999 7625 12025 7631
rect 8751 7601 8777 7607
rect 11047 7601 11073 7607
rect 8409 7575 8415 7601
rect 8441 7575 8447 7601
rect 10817 7575 10823 7601
rect 10849 7575 10855 7601
rect 8751 7569 8777 7575
rect 11047 7569 11073 7575
rect 11775 7601 11801 7607
rect 14065 7575 14071 7601
rect 14097 7575 14103 7601
rect 11775 7569 11801 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9311 7321 9337 7327
rect 13007 7321 13033 7327
rect 8017 7295 8023 7321
rect 8049 7295 8055 7321
rect 9081 7295 9087 7321
rect 9113 7295 9119 7321
rect 11713 7295 11719 7321
rect 11745 7295 11751 7321
rect 12777 7295 12783 7321
rect 12809 7295 12815 7321
rect 9311 7289 9337 7295
rect 13007 7289 13033 7295
rect 10879 7265 10905 7271
rect 7681 7239 7687 7265
rect 7713 7239 7719 7265
rect 11377 7239 11383 7265
rect 11409 7239 11415 7265
rect 10879 7233 10905 7239
rect 10711 7209 10737 7215
rect 10711 7177 10737 7183
rect 10767 7153 10793 7159
rect 10767 7121 10793 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 11551 6985 11577 6991
rect 11551 6953 11577 6959
rect 10929 6903 10935 6929
rect 10961 6903 10967 6929
rect 11321 6847 11327 6873
rect 11353 6847 11359 6873
rect 9865 6791 9871 6817
rect 9897 6791 9903 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8857 2143 8863 2169
rect 8889 2143 8895 2169
rect 10537 2143 10543 2169
rect 10569 2143 10575 2169
rect 9367 2057 9393 2063
rect 9367 2025 9393 2031
rect 11047 2057 11073 2063
rect 11047 2025 11073 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 13063 1833 13089 1839
rect 13063 1801 13089 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10705 1751 10711 1777
rect 10737 1751 10743 1777
rect 12609 1751 12615 1777
rect 12641 1751 12647 1777
rect 11215 1665 11241 1671
rect 11215 1633 11241 1639
rect 17263 1665 17289 1671
rect 17263 1633 17289 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9591 19111 9617 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 9871 18999 9897 19025
rect 10711 18999 10737 19025
rect 12279 18999 12305 19025
rect 13735 18943 13761 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9367 18719 9393 18745
rect 11047 18719 11073 18745
rect 13119 18719 13145 18745
rect 8863 18607 8889 18633
rect 10655 18607 10681 18633
rect 12615 18607 12641 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 13399 18327 13425 18353
rect 12895 18215 12921 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9927 14407 9953 14433
rect 11663 14407 11689 14433
rect 12223 14295 12249 14321
rect 9983 14239 10009 14265
rect 10207 14239 10233 14265
rect 10263 14239 10289 14265
rect 11607 14239 11633 14265
rect 12335 14239 12361 14265
rect 9927 14183 9953 14209
rect 10095 14183 10121 14209
rect 11663 14183 11689 14209
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 12671 14015 12697 14041
rect 9591 13959 9617 13985
rect 11271 13959 11297 13985
rect 9255 13903 9281 13929
rect 10879 13903 10905 13929
rect 12615 13903 12641 13929
rect 13007 13903 13033 13929
rect 10655 13847 10681 13873
rect 12335 13847 12361 13873
rect 12671 13791 12697 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9983 13567 10009 13593
rect 10767 13567 10793 13593
rect 12895 13567 12921 13593
rect 13119 13567 13145 13593
rect 8359 13511 8385 13537
rect 8527 13511 8553 13537
rect 10151 13511 10177 13537
rect 11439 13511 11465 13537
rect 8919 13455 8945 13481
rect 10263 13455 10289 13481
rect 10319 13455 10345 13481
rect 11831 13455 11857 13481
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 9143 13231 9169 13257
rect 10319 13231 10345 13257
rect 11551 13231 11577 13257
rect 11663 13231 11689 13257
rect 11831 13231 11857 13257
rect 8751 13175 8777 13201
rect 9255 13175 9281 13201
rect 9311 13175 9337 13201
rect 11719 13175 11745 13201
rect 11943 13175 11969 13201
rect 11999 13175 12025 13201
rect 7015 13119 7041 13145
rect 10151 13119 10177 13145
rect 18831 13119 18857 13145
rect 7351 13063 7377 13089
rect 8415 13063 8441 13089
rect 19951 13063 19977 13089
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 967 12783 993 12809
rect 4999 12783 5025 12809
rect 8527 12783 8553 12809
rect 20007 12783 20033 12809
rect 2143 12727 2169 12753
rect 6455 12727 6481 12753
rect 8639 12727 8665 12753
rect 12783 12727 12809 12753
rect 12951 12727 12977 12753
rect 18831 12727 18857 12753
rect 6063 12671 6089 12697
rect 6791 12671 6817 12697
rect 7967 12671 7993 12697
rect 8135 12671 8161 12697
rect 10655 12671 10681 12697
rect 13007 12671 13033 12697
rect 6735 12615 6761 12641
rect 7015 12615 7041 12641
rect 8807 12615 8833 12641
rect 10711 12615 10737 12641
rect 10823 12615 10849 12641
rect 12615 12615 12641 12641
rect 12727 12615 12753 12641
rect 13119 12615 13145 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8695 12447 8721 12473
rect 12223 12447 12249 12473
rect 6567 12391 6593 12417
rect 14407 12391 14433 12417
rect 2143 12335 2169 12361
rect 6959 12335 6985 12361
rect 9031 12335 9057 12361
rect 11271 12335 11297 12361
rect 12055 12335 12081 12361
rect 12111 12335 12137 12361
rect 12335 12335 12361 12361
rect 12671 12335 12697 12361
rect 14295 12335 14321 12361
rect 18831 12335 18857 12361
rect 5503 12279 5529 12305
rect 7183 12279 7209 12305
rect 9143 12279 9169 12305
rect 9815 12279 9841 12305
rect 10879 12279 10905 12305
rect 11495 12279 11521 12305
rect 12391 12279 12417 12305
rect 13007 12279 13033 12305
rect 14071 12279 14097 12305
rect 14631 12279 14657 12305
rect 967 12223 993 12249
rect 8919 12223 8945 12249
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 6399 12055 6425 12081
rect 967 11999 993 12025
rect 6903 11999 6929 12025
rect 7575 11999 7601 12025
rect 10879 11999 10905 12025
rect 13399 11999 13425 12025
rect 2143 11943 2169 11969
rect 6455 11943 6481 11969
rect 6959 11943 6985 11969
rect 9031 11943 9057 11969
rect 9143 11943 9169 11969
rect 9311 11943 9337 11969
rect 10655 11943 10681 11969
rect 11663 11943 11689 11969
rect 11999 11943 12025 11969
rect 13623 11943 13649 11969
rect 7183 11887 7209 11913
rect 8639 11887 8665 11913
rect 9255 11887 9281 11913
rect 9479 11887 9505 11913
rect 11551 11887 11577 11913
rect 12335 11887 12361 11913
rect 6903 11831 6929 11857
rect 7071 11831 7097 11857
rect 9703 11831 9729 11857
rect 10767 11831 10793 11857
rect 10879 11831 10905 11857
rect 11775 11831 11801 11857
rect 11831 11831 11857 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 6959 11663 6985 11689
rect 8807 11663 8833 11689
rect 8863 11663 8889 11689
rect 9367 11663 9393 11689
rect 10375 11663 10401 11689
rect 11719 11663 11745 11689
rect 11999 11663 12025 11689
rect 9255 11607 9281 11633
rect 9927 11607 9953 11633
rect 6847 11551 6873 11577
rect 6903 11551 6929 11577
rect 7015 11551 7041 11577
rect 7071 11551 7097 11577
rect 8751 11551 8777 11577
rect 8919 11551 8945 11577
rect 9031 11551 9057 11577
rect 9199 11551 9225 11577
rect 9871 11551 9897 11577
rect 10039 11551 10065 11577
rect 10487 11551 10513 11577
rect 11887 11551 11913 11577
rect 12111 11551 12137 11577
rect 12223 11551 12249 11577
rect 10319 11495 10345 11521
rect 11439 11495 11465 11521
rect 11551 11495 11577 11521
rect 12279 11495 12305 11521
rect 12671 11495 12697 11521
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 12559 11271 12585 11297
rect 967 11215 993 11241
rect 14239 11215 14265 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 6735 11159 6761 11185
rect 6959 11159 6985 11185
rect 7183 11159 7209 11185
rect 7351 11159 7377 11185
rect 7967 11159 7993 11185
rect 8247 11159 8273 11185
rect 8919 11159 8945 11185
rect 9143 11159 9169 11185
rect 9591 11159 9617 11185
rect 9815 11159 9841 11185
rect 10263 11159 10289 11185
rect 11047 11159 11073 11185
rect 12279 11159 12305 11185
rect 12503 11159 12529 11185
rect 12783 11159 12809 11185
rect 18831 11159 18857 11185
rect 6903 11103 6929 11129
rect 9479 11103 9505 11129
rect 10319 11103 10345 11129
rect 11215 11103 11241 11129
rect 12615 11103 12641 11129
rect 13175 11103 13201 11129
rect 6791 11047 6817 11073
rect 7239 11047 7265 11073
rect 8079 11047 8105 11073
rect 8303 11047 8329 11073
rect 8751 11047 8777 11073
rect 8975 11047 9001 11073
rect 9871 11047 9897 11073
rect 11159 11047 11185 11073
rect 12391 11047 12417 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 11887 10879 11913 10905
rect 12279 10879 12305 10905
rect 12671 10879 12697 10905
rect 13119 10879 13145 10905
rect 13231 10879 13257 10905
rect 8863 10823 8889 10849
rect 6343 10767 6369 10793
rect 8415 10767 8441 10793
rect 8751 10767 8777 10793
rect 9255 10767 9281 10793
rect 11999 10767 12025 10793
rect 12223 10767 12249 10793
rect 12391 10767 12417 10793
rect 12783 10767 12809 10793
rect 12895 10767 12921 10793
rect 13063 10767 13089 10793
rect 6679 10711 6705 10737
rect 7743 10711 7769 10737
rect 7967 10711 7993 10737
rect 8191 10711 8217 10737
rect 10823 10711 10849 10737
rect 12839 10711 12865 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 4999 10431 5025 10457
rect 6063 10431 6089 10457
rect 6791 10431 6817 10457
rect 7967 10431 7993 10457
rect 10039 10431 10065 10457
rect 6455 10375 6481 10401
rect 9815 10375 9841 10401
rect 10207 10375 10233 10401
rect 10823 10375 10849 10401
rect 12839 10319 12865 10345
rect 9983 10263 10009 10289
rect 10095 10263 10121 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 6791 10039 6817 10065
rect 6959 10039 6985 10065
rect 7071 10039 7097 10065
rect 7351 10039 7377 10065
rect 8695 10039 8721 10065
rect 10375 10039 10401 10065
rect 10711 10039 10737 10065
rect 11103 10039 11129 10065
rect 11439 10039 11465 10065
rect 11607 10039 11633 10065
rect 11775 10039 11801 10065
rect 13847 10039 13873 10065
rect 6903 9983 6929 10009
rect 7015 9983 7041 10009
rect 7799 9983 7825 10009
rect 8863 9983 8889 10009
rect 9087 9983 9113 10009
rect 9255 9983 9281 10009
rect 9983 9983 10009 10009
rect 10263 9983 10289 10009
rect 10543 9983 10569 10009
rect 10879 9983 10905 10009
rect 10991 9983 11017 10009
rect 11271 9983 11297 10009
rect 12335 9983 12361 10009
rect 14183 9983 14209 10009
rect 6511 9927 6537 9953
rect 7295 9927 7321 9953
rect 7463 9927 7489 9953
rect 7911 9927 7937 9953
rect 8135 9927 8161 9953
rect 8751 9927 8777 9953
rect 9759 9927 9785 9953
rect 10935 9927 10961 9953
rect 12783 9927 12809 9953
rect 9087 9871 9113 9897
rect 12167 9871 12193 9897
rect 12335 9871 12361 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 7015 9703 7041 9729
rect 11047 9703 11073 9729
rect 11439 9703 11465 9729
rect 5335 9647 5361 9673
rect 6399 9647 6425 9673
rect 7183 9647 7209 9673
rect 8807 9647 8833 9673
rect 11215 9647 11241 9673
rect 12055 9647 12081 9673
rect 13231 9647 13257 9673
rect 14295 9647 14321 9673
rect 20007 9647 20033 9673
rect 4999 9591 5025 9617
rect 6735 9591 6761 9617
rect 6847 9591 6873 9617
rect 8023 9591 8049 9617
rect 8471 9591 8497 9617
rect 8695 9591 8721 9617
rect 8919 9591 8945 9617
rect 9031 9591 9057 9617
rect 9367 9591 9393 9617
rect 9703 9591 9729 9617
rect 9927 9591 9953 9617
rect 10319 9591 10345 9617
rect 10767 9591 10793 9617
rect 11999 9591 12025 9617
rect 12335 9591 12361 9617
rect 12839 9591 12865 9617
rect 18831 9591 18857 9617
rect 7239 9535 7265 9561
rect 8079 9535 8105 9561
rect 8303 9535 8329 9561
rect 9647 9535 9673 9561
rect 10375 9535 10401 9561
rect 11159 9535 11185 9561
rect 11383 9535 11409 9561
rect 11775 9535 11801 9561
rect 12447 9535 12473 9561
rect 8191 9479 8217 9505
rect 9255 9479 9281 9505
rect 10823 9479 10849 9505
rect 10935 9479 10961 9505
rect 11439 9479 11465 9505
rect 11887 9479 11913 9505
rect 12055 9479 12081 9505
rect 12671 9479 12697 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 6287 9311 6313 9337
rect 7183 9311 7209 9337
rect 8359 9311 8385 9337
rect 9143 9311 9169 9337
rect 9591 9311 9617 9337
rect 10431 9311 10457 9337
rect 11327 9311 11353 9337
rect 13007 9311 13033 9337
rect 8415 9255 8441 9281
rect 8695 9255 8721 9281
rect 9535 9255 9561 9281
rect 10151 9255 10177 9281
rect 10823 9255 10849 9281
rect 10879 9255 10905 9281
rect 11495 9255 11521 9281
rect 12615 9255 12641 9281
rect 6455 9199 6481 9225
rect 6567 9199 6593 9225
rect 7015 9199 7041 9225
rect 8807 9199 8833 9225
rect 8975 9199 9001 9225
rect 9087 9199 9113 9225
rect 9367 9199 9393 9225
rect 9759 9199 9785 9225
rect 9871 9199 9897 9225
rect 10319 9199 10345 9225
rect 12727 9199 12753 9225
rect 12895 9199 12921 9225
rect 13231 9199 13257 9225
rect 13343 9199 13369 9225
rect 18943 9199 18969 9225
rect 6007 9143 6033 9169
rect 9311 9143 9337 9169
rect 10487 9143 10513 9169
rect 12335 9143 12361 9169
rect 6791 9087 6817 9113
rect 8359 9087 8385 9113
rect 10879 9087 10905 9113
rect 12895 9087 12921 9113
rect 13175 9087 13201 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 6063 8919 6089 8945
rect 11047 8919 11073 8945
rect 6119 8863 6145 8889
rect 7015 8863 7041 8889
rect 13231 8863 13257 8889
rect 14295 8863 14321 8889
rect 20007 8863 20033 8889
rect 6903 8807 6929 8833
rect 7295 8807 7321 8833
rect 9927 8807 9953 8833
rect 10991 8807 11017 8833
rect 12839 8807 12865 8833
rect 14631 8807 14657 8833
rect 18831 8807 18857 8833
rect 6287 8751 6313 8777
rect 9983 8751 10009 8777
rect 10767 8751 10793 8777
rect 6455 8695 6481 8721
rect 10095 8695 10121 8721
rect 10599 8695 10625 8721
rect 10711 8695 10737 8721
rect 11047 8695 11073 8721
rect 12671 8695 12697 8721
rect 14743 8695 14769 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 8303 8527 8329 8553
rect 8975 8527 9001 8553
rect 9759 8527 9785 8553
rect 10151 8527 10177 8553
rect 10207 8527 10233 8553
rect 5839 8471 5865 8497
rect 7463 8471 7489 8497
rect 7631 8471 7657 8497
rect 8079 8471 8105 8497
rect 8919 8471 8945 8497
rect 9591 8471 9617 8497
rect 11607 8471 11633 8497
rect 11887 8471 11913 8497
rect 5503 8415 5529 8441
rect 8191 8415 8217 8441
rect 8695 8415 8721 8441
rect 9087 8415 9113 8441
rect 10319 8415 10345 8441
rect 10431 8415 10457 8441
rect 11663 8415 11689 8441
rect 11775 8415 11801 8441
rect 6903 8359 6929 8385
rect 7127 8359 7153 8385
rect 8919 8359 8945 8385
rect 10263 8359 10289 8385
rect 8135 8303 8161 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 12727 8135 12753 8161
rect 20007 8079 20033 8105
rect 8303 8023 8329 8049
rect 8415 8023 8441 8049
rect 8639 8023 8665 8049
rect 10599 8023 10625 8049
rect 12167 8023 12193 8049
rect 12279 8023 12305 8049
rect 12391 8023 12417 8049
rect 12447 8023 12473 8049
rect 12783 8023 12809 8049
rect 18831 8023 18857 8049
rect 10711 7967 10737 7993
rect 10767 7967 10793 7993
rect 8359 7911 8385 7937
rect 10991 7911 11017 7937
rect 12559 7911 12585 7937
rect 12839 7911 12865 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8863 7743 8889 7769
rect 9031 7743 9057 7769
rect 12167 7743 12193 7769
rect 14295 7743 14321 7769
rect 7351 7687 7377 7713
rect 8919 7687 8945 7713
rect 9759 7687 9785 7713
rect 11159 7687 11185 7713
rect 11271 7687 11297 7713
rect 11887 7687 11913 7713
rect 12279 7687 12305 7713
rect 12335 7687 12361 7713
rect 13007 7687 13033 7713
rect 7015 7631 7041 7657
rect 9199 7631 9225 7657
rect 9423 7631 9449 7657
rect 10935 7631 10961 7657
rect 11663 7631 11689 7657
rect 11999 7631 12025 7657
rect 12615 7631 12641 7657
rect 8415 7575 8441 7601
rect 8751 7575 8777 7601
rect 10823 7575 10849 7601
rect 11047 7575 11073 7601
rect 11775 7575 11801 7601
rect 14071 7575 14097 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8023 7295 8049 7321
rect 9087 7295 9113 7321
rect 9311 7295 9337 7321
rect 11719 7295 11745 7321
rect 12783 7295 12809 7321
rect 13007 7295 13033 7321
rect 7687 7239 7713 7265
rect 10879 7239 10905 7265
rect 11383 7239 11409 7265
rect 10711 7183 10737 7209
rect 10767 7127 10793 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 11551 6959 11577 6985
rect 10935 6903 10961 6929
rect 11327 6847 11353 6873
rect 9871 6791 9897 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8863 2143 8889 2169
rect 10543 2143 10569 2169
rect 9367 2031 9393 2057
rect 11047 2031 11073 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 13063 1807 13089 1833
rect 8807 1751 8833 1777
rect 10711 1751 10737 1777
rect 12615 1751 12641 1777
rect 11215 1639 11241 1665
rect 17263 1639 17289 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8736 20600 8792 21000
rect 9744 20600 9800 21000
rect 10416 20600 10472 21000
rect 11088 20600 11144 21000
rect 12096 20600 12152 21000
rect 12432 20600 12488 21000
rect 12768 20600 12824 21000
rect 13104 20600 13160 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8750 18746 8778 20600
rect 9758 19334 9786 20600
rect 9590 19306 9786 19334
rect 9590 19137 9618 19306
rect 9590 19111 9591 19137
rect 9617 19111 9618 19137
rect 9590 19105 9618 19111
rect 9870 19026 9898 19031
rect 9814 19025 9898 19026
rect 9814 18999 9871 19025
rect 9897 18999 9898 19025
rect 9814 18998 9898 18999
rect 8750 18713 8778 18718
rect 9366 18746 9394 18751
rect 9366 18699 9394 18718
rect 8862 18634 8890 18639
rect 8414 18633 8890 18634
rect 8414 18607 8863 18633
rect 8889 18607 8890 18633
rect 8414 18606 8890 18607
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2086 13818 2114 13823
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11241 994 11247
rect 966 11215 967 11241
rect 993 11215 994 11241
rect 966 10794 994 11215
rect 2086 11074 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8358 13538 8386 13543
rect 8358 13491 8386 13510
rect 7014 13145 7042 13151
rect 7014 13119 7015 13145
rect 7041 13119 7042 13145
rect 7014 13090 7042 13119
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 4998 12810 5026 12815
rect 4998 12763 5026 12782
rect 6902 12810 6930 12815
rect 2142 12754 2170 12759
rect 2142 12707 2170 12726
rect 6454 12753 6482 12759
rect 6454 12727 6455 12753
rect 6481 12727 6482 12753
rect 6062 12698 6090 12703
rect 6062 12697 6426 12698
rect 6062 12671 6063 12697
rect 6089 12671 6426 12697
rect 6062 12670 6426 12671
rect 6062 12665 6090 12670
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 5502 12306 5530 12311
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 5502 12082 5530 12278
rect 5502 12049 5530 12054
rect 6398 12081 6426 12670
rect 6454 12642 6482 12727
rect 6790 12698 6818 12703
rect 6790 12697 6874 12698
rect 6790 12671 6791 12697
rect 6817 12671 6874 12697
rect 6790 12670 6874 12671
rect 6790 12665 6818 12670
rect 6734 12642 6762 12647
rect 6454 12609 6482 12614
rect 6566 12641 6762 12642
rect 6566 12615 6735 12641
rect 6761 12615 6762 12641
rect 6566 12614 6762 12615
rect 6566 12417 6594 12614
rect 6734 12609 6762 12614
rect 6566 12391 6567 12417
rect 6593 12391 6594 12417
rect 6566 12385 6594 12391
rect 6398 12055 6399 12081
rect 6425 12055 6426 12081
rect 6398 12049 6426 12055
rect 6790 12082 6818 12087
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 6454 11970 6482 11975
rect 6454 11923 6482 11942
rect 6790 11466 6818 12054
rect 6846 11690 6874 12670
rect 6902 12250 6930 12782
rect 7014 12642 7042 13062
rect 7350 13089 7378 13095
rect 7350 13063 7351 13089
rect 7377 13063 7378 13089
rect 7350 12698 7378 13063
rect 8414 13090 8442 18606
rect 8862 18601 8890 18606
rect 9590 14434 9618 14439
rect 9310 14210 9338 14215
rect 9254 13930 9282 13935
rect 9254 13883 9282 13902
rect 8526 13538 8554 13543
rect 8526 13454 8554 13510
rect 8918 13481 8946 13487
rect 8918 13455 8919 13481
rect 8945 13455 8946 13481
rect 8918 13454 8946 13455
rect 8526 13426 8610 13454
rect 8918 13426 9170 13454
rect 8582 13202 8610 13426
rect 9142 13257 9170 13426
rect 9142 13231 9143 13257
rect 9169 13231 9170 13257
rect 9142 13225 9170 13231
rect 8750 13202 8778 13207
rect 8582 13201 8778 13202
rect 8582 13175 8751 13201
rect 8777 13175 8778 13201
rect 8582 13174 8778 13175
rect 8582 13090 8610 13174
rect 8750 13169 8778 13174
rect 9254 13201 9282 13207
rect 9254 13175 9255 13201
rect 9281 13175 9282 13201
rect 8414 13089 8554 13090
rect 8414 13063 8415 13089
rect 8441 13063 8554 13089
rect 8414 13062 8554 13063
rect 8414 13057 8442 13062
rect 8526 12809 8554 13062
rect 8582 13057 8610 13062
rect 8526 12783 8527 12809
rect 8553 12783 8554 12809
rect 8526 12777 8554 12783
rect 8638 12754 8666 12759
rect 8638 12707 8666 12726
rect 7350 12665 7378 12670
rect 7966 12698 7994 12703
rect 7966 12651 7994 12670
rect 8134 12697 8162 12703
rect 8134 12671 8135 12697
rect 8161 12671 8162 12697
rect 6958 12361 6986 12367
rect 6958 12335 6959 12361
rect 6985 12335 6986 12361
rect 6958 12306 6986 12335
rect 7014 12306 7042 12614
rect 8134 12474 8162 12671
rect 8806 12642 8834 12647
rect 8806 12641 9058 12642
rect 8806 12615 8807 12641
rect 8833 12615 9058 12641
rect 8806 12614 9058 12615
rect 8806 12609 8834 12614
rect 8134 12441 8162 12446
rect 8694 12474 8722 12479
rect 8694 12427 8722 12446
rect 9030 12361 9058 12614
rect 9030 12335 9031 12361
rect 9057 12335 9058 12361
rect 9030 12329 9058 12335
rect 7182 12306 7210 12311
rect 6958 12305 7210 12306
rect 6958 12279 7183 12305
rect 7209 12279 7210 12305
rect 6958 12278 7210 12279
rect 6902 12222 6986 12250
rect 6902 12025 6930 12031
rect 6902 11999 6903 12025
rect 6929 11999 6930 12025
rect 6902 11970 6930 11999
rect 6902 11937 6930 11942
rect 6958 11969 6986 12222
rect 6958 11943 6959 11969
rect 6985 11943 6986 11969
rect 6958 11937 6986 11943
rect 6902 11857 6930 11863
rect 6902 11831 6903 11857
rect 6929 11831 6930 11857
rect 6902 11802 6930 11831
rect 6902 11769 6930 11774
rect 7070 11857 7098 11863
rect 7070 11831 7071 11857
rect 7097 11831 7098 11857
rect 6958 11690 6986 11695
rect 7070 11690 7098 11831
rect 7126 11802 7154 12278
rect 7182 12273 7210 12278
rect 9142 12306 9170 12311
rect 9142 12305 9226 12306
rect 9142 12279 9143 12305
rect 9169 12279 9226 12305
rect 9142 12278 9226 12279
rect 9142 12273 9170 12278
rect 8918 12250 8946 12255
rect 8582 12249 8946 12250
rect 8582 12223 8919 12249
rect 8945 12223 8946 12249
rect 8582 12222 8946 12223
rect 7574 12026 7602 12031
rect 7574 11979 7602 11998
rect 7182 11914 7210 11919
rect 7182 11913 7434 11914
rect 7182 11887 7183 11913
rect 7209 11887 7434 11913
rect 7182 11886 7434 11887
rect 7182 11881 7210 11886
rect 7126 11774 7322 11802
rect 6846 11689 6986 11690
rect 6846 11663 6959 11689
rect 6985 11663 6986 11689
rect 6846 11662 6986 11663
rect 6958 11657 6986 11662
rect 7014 11662 7098 11690
rect 6846 11578 6874 11583
rect 6846 11531 6874 11550
rect 6902 11577 6930 11583
rect 6902 11551 6903 11577
rect 6929 11551 6930 11577
rect 6902 11466 6930 11551
rect 7014 11577 7042 11662
rect 7014 11551 7015 11577
rect 7041 11551 7042 11577
rect 7014 11522 7042 11551
rect 7014 11489 7042 11494
rect 7070 11577 7098 11583
rect 7070 11551 7071 11577
rect 7097 11551 7098 11577
rect 6790 11438 6930 11466
rect 6734 11410 6762 11415
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 4998 11186 5026 11191
rect 2086 11041 2114 11046
rect 966 10761 994 10766
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 4998 10457 5026 11158
rect 6734 11185 6762 11382
rect 7014 11410 7042 11415
rect 6734 11159 6735 11185
rect 6761 11159 6762 11185
rect 6734 11153 6762 11159
rect 6958 11185 6986 11191
rect 6958 11159 6959 11185
rect 6985 11159 6986 11185
rect 6902 11130 6930 11135
rect 6902 11083 6930 11102
rect 6790 11073 6818 11079
rect 6790 11047 6791 11073
rect 6817 11047 6818 11073
rect 4998 10431 4999 10457
rect 5025 10431 5026 10457
rect 4998 10402 5026 10431
rect 6062 10962 6090 10967
rect 6062 10457 6090 10934
rect 6790 10962 6818 11047
rect 6790 10929 6818 10934
rect 6062 10431 6063 10457
rect 6089 10431 6090 10457
rect 6062 10425 6090 10431
rect 6342 10793 6370 10799
rect 6342 10767 6343 10793
rect 6369 10767 6370 10793
rect 6342 10458 6370 10767
rect 6678 10737 6706 10743
rect 6678 10711 6679 10737
rect 6705 10711 6706 10737
rect 6454 10458 6482 10463
rect 6342 10430 6454 10458
rect 4998 10369 5026 10374
rect 6454 10401 6482 10430
rect 6454 10375 6455 10401
rect 6481 10375 6482 10401
rect 6454 10094 6482 10375
rect 6454 10066 6538 10094
rect 6510 9953 6538 10066
rect 6510 9927 6511 9953
rect 6537 9927 6538 9953
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 5334 9674 5362 9679
rect 5334 9627 5362 9646
rect 6398 9673 6426 9679
rect 6398 9647 6399 9673
rect 6425 9647 6426 9673
rect 4998 9617 5026 9623
rect 6398 9618 6426 9647
rect 4998 9591 4999 9617
rect 5025 9591 5026 9617
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 4998 8442 5026 9591
rect 6286 9590 6398 9618
rect 6286 9337 6314 9590
rect 6398 9585 6426 9590
rect 6286 9311 6287 9337
rect 6313 9311 6314 9337
rect 6286 9305 6314 9311
rect 6062 9226 6090 9231
rect 6006 9170 6034 9175
rect 6006 9123 6034 9142
rect 6062 8946 6090 9198
rect 6454 9225 6482 9231
rect 6454 9199 6455 9225
rect 6481 9199 6482 9225
rect 6454 9170 6482 9199
rect 6454 9137 6482 9142
rect 5838 8945 6090 8946
rect 5838 8919 6063 8945
rect 6089 8919 6090 8945
rect 5838 8918 6090 8919
rect 5838 8497 5866 8918
rect 6062 8913 6090 8918
rect 6286 9114 6314 9119
rect 6118 8890 6146 8895
rect 6286 8890 6314 9086
rect 6118 8889 6314 8890
rect 6118 8863 6119 8889
rect 6145 8863 6314 8889
rect 6118 8862 6314 8863
rect 6118 8857 6146 8862
rect 6286 8777 6314 8862
rect 6286 8751 6287 8777
rect 6313 8751 6314 8777
rect 6286 8745 6314 8751
rect 5838 8471 5839 8497
rect 5865 8471 5866 8497
rect 5838 8465 5866 8471
rect 6454 8721 6482 8727
rect 6454 8695 6455 8721
rect 6481 8695 6482 8721
rect 6454 8498 6482 8695
rect 6454 8465 6482 8470
rect 4998 8409 5026 8414
rect 5502 8442 5530 8447
rect 5502 8395 5530 8414
rect 6510 8442 6538 9927
rect 6678 9954 6706 10711
rect 6790 10458 6818 10463
rect 6790 10411 6818 10430
rect 6734 10402 6762 10407
rect 6734 10094 6762 10374
rect 6734 10066 6818 10094
rect 6790 10065 6818 10066
rect 6790 10039 6791 10065
rect 6817 10039 6818 10065
rect 6790 10033 6818 10039
rect 6846 10066 6874 10071
rect 6678 9921 6706 9926
rect 6846 9730 6874 10038
rect 6958 10065 6986 11159
rect 6958 10039 6959 10065
rect 6985 10039 6986 10065
rect 6958 10033 6986 10039
rect 6902 10009 6930 10015
rect 6902 9983 6903 10009
rect 6929 9983 6930 10009
rect 6902 9898 6930 9983
rect 7014 10010 7042 11382
rect 7070 10066 7098 11551
rect 7182 11522 7210 11527
rect 7182 11242 7210 11494
rect 7182 11185 7210 11214
rect 7182 11159 7183 11185
rect 7209 11159 7210 11185
rect 7182 11153 7210 11159
rect 7070 10019 7098 10038
rect 7126 11130 7154 11135
rect 7014 9963 7042 9982
rect 7126 9954 7154 11102
rect 7238 11073 7266 11079
rect 7238 11047 7239 11073
rect 7265 11047 7266 11073
rect 7238 10094 7266 11047
rect 7294 10458 7322 11774
rect 7350 11186 7378 11191
rect 7350 11139 7378 11158
rect 7406 10794 7434 11886
rect 7966 11186 7994 11191
rect 8246 11186 8274 11191
rect 7406 10761 7434 10766
rect 7742 11185 8274 11186
rect 7742 11159 7967 11185
rect 7993 11159 8247 11185
rect 8273 11159 8274 11185
rect 7742 11158 8274 11159
rect 7742 10737 7770 11158
rect 7966 11153 7994 11158
rect 8246 11153 8274 11158
rect 8078 11073 8106 11079
rect 8078 11047 8079 11073
rect 8105 11047 8106 11073
rect 7742 10711 7743 10737
rect 7769 10711 7770 10737
rect 7742 10705 7770 10711
rect 7798 10962 7826 10967
rect 7294 10425 7322 10430
rect 6902 9865 6930 9870
rect 7070 9926 7154 9954
rect 7182 10066 7266 10094
rect 6790 9702 6874 9730
rect 7014 9730 7042 9735
rect 6734 9617 6762 9623
rect 6734 9591 6735 9617
rect 6761 9591 6762 9617
rect 6566 9226 6594 9231
rect 6566 9179 6594 9198
rect 6734 9114 6762 9591
rect 6734 9081 6762 9086
rect 6790 9113 6818 9702
rect 7014 9683 7042 9702
rect 6846 9618 6874 9623
rect 6846 9226 6874 9590
rect 7070 9394 7098 9926
rect 7182 9674 7210 10066
rect 7350 10065 7378 10071
rect 7350 10039 7351 10065
rect 7377 10039 7378 10065
rect 7350 10010 7378 10039
rect 7294 9954 7322 9959
rect 7294 9907 7322 9926
rect 7182 9627 7210 9646
rect 7238 9562 7266 9567
rect 7350 9562 7378 9982
rect 7406 10066 7434 10071
rect 7406 9618 7434 10038
rect 7798 10009 7826 10934
rect 7966 10737 7994 10743
rect 7966 10711 7967 10737
rect 7993 10711 7994 10737
rect 7798 9983 7799 10009
rect 7825 9983 7826 10009
rect 7798 9977 7826 9983
rect 7910 10570 7938 10575
rect 7462 9954 7490 9959
rect 7462 9907 7490 9926
rect 7910 9953 7938 10542
rect 7966 10458 7994 10711
rect 7966 10411 7994 10430
rect 8078 10066 8106 11047
rect 8302 11073 8330 11079
rect 8302 11047 8303 11073
rect 8329 11047 8330 11073
rect 8190 10962 8218 10967
rect 8190 10737 8218 10934
rect 8302 10794 8330 11047
rect 8414 10794 8442 10799
rect 8302 10766 8414 10794
rect 8414 10747 8442 10766
rect 8190 10711 8191 10737
rect 8217 10711 8218 10737
rect 8190 10705 8218 10711
rect 8582 10178 8610 12222
rect 8918 12217 8946 12222
rect 8806 12026 8834 12031
rect 8638 11914 8666 11919
rect 8638 11867 8666 11886
rect 8694 11746 8722 11751
rect 8694 11018 8722 11718
rect 8806 11689 8834 11998
rect 9030 11969 9058 11975
rect 9030 11943 9031 11969
rect 9057 11943 9058 11969
rect 9030 11858 9058 11943
rect 9030 11825 9058 11830
rect 9142 11969 9170 11975
rect 9142 11943 9143 11969
rect 9169 11943 9170 11969
rect 8806 11663 8807 11689
rect 8833 11663 8834 11689
rect 8806 11657 8834 11663
rect 8862 11690 8890 11695
rect 9142 11690 9170 11943
rect 9198 11970 9226 12278
rect 9254 12194 9282 13175
rect 9310 13201 9338 14182
rect 9590 13985 9618 14406
rect 9814 14322 9842 18998
rect 9870 18993 9898 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10430 18746 10458 20600
rect 11102 19334 11130 20600
rect 11102 19306 11242 19334
rect 11214 19137 11242 19306
rect 11214 19111 11215 19137
rect 11241 19111 11242 19137
rect 11214 19105 11242 19111
rect 12110 19138 12138 20600
rect 12110 19105 12138 19110
rect 10430 18713 10458 18718
rect 10710 19025 10738 19031
rect 12278 19026 12306 19031
rect 10710 18999 10711 19025
rect 10737 18999 10738 19025
rect 10654 18633 10682 18639
rect 10654 18607 10655 18633
rect 10681 18607 10682 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9926 14434 9954 14439
rect 9926 14387 9954 14406
rect 9814 14289 9842 14294
rect 10038 14294 10178 14322
rect 9982 14266 10010 14271
rect 10038 14266 10066 14294
rect 9982 14265 10066 14266
rect 9982 14239 9983 14265
rect 10009 14239 10066 14265
rect 9982 14238 10066 14239
rect 9982 14233 10010 14238
rect 9926 14210 9954 14215
rect 9590 13959 9591 13985
rect 9617 13959 9618 13985
rect 9590 13953 9618 13959
rect 9814 14209 9954 14210
rect 9814 14183 9927 14209
rect 9953 14183 9954 14209
rect 9814 14182 9954 14183
rect 9310 13175 9311 13201
rect 9337 13175 9338 13201
rect 9310 13169 9338 13175
rect 9814 12978 9842 14182
rect 9926 14177 9954 14182
rect 10094 14210 10122 14215
rect 10094 14163 10122 14182
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9982 14042 10010 14047
rect 9982 13593 10010 14014
rect 9982 13567 9983 13593
rect 10009 13567 10010 13593
rect 9982 13561 10010 13567
rect 10150 13537 10178 14294
rect 10206 14266 10234 14271
rect 10206 14042 10234 14238
rect 10206 14009 10234 14014
rect 10262 14265 10290 14271
rect 10262 14239 10263 14265
rect 10289 14239 10290 14265
rect 10262 13874 10290 14239
rect 10654 13874 10682 18607
rect 10150 13511 10151 13537
rect 10177 13511 10178 13537
rect 10150 13505 10178 13511
rect 10206 13846 10290 13874
rect 10318 13873 10682 13874
rect 10318 13847 10655 13873
rect 10681 13847 10682 13873
rect 10318 13846 10682 13847
rect 10206 13370 10234 13846
rect 10318 13818 10346 13846
rect 10654 13841 10682 13846
rect 10262 13790 10346 13818
rect 10262 13481 10290 13790
rect 10262 13455 10263 13481
rect 10289 13455 10290 13481
rect 10262 13449 10290 13455
rect 10318 13481 10346 13487
rect 10318 13455 10319 13481
rect 10345 13455 10346 13481
rect 10318 13370 10346 13455
rect 9918 13342 10050 13347
rect 10206 13342 10346 13370
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10318 13258 10346 13342
rect 10318 13211 10346 13230
rect 9758 12950 9842 12978
rect 10150 13145 10178 13151
rect 10150 13119 10151 13145
rect 10177 13119 10178 13145
rect 9422 12754 9450 12759
rect 9254 12166 9338 12194
rect 9198 11937 9226 11942
rect 9310 11969 9338 12166
rect 9310 11943 9311 11969
rect 9337 11943 9338 11969
rect 9254 11914 9282 11919
rect 9254 11867 9282 11886
rect 8862 11689 9170 11690
rect 8862 11663 8863 11689
rect 8889 11663 9170 11689
rect 8862 11662 9170 11663
rect 9310 11690 9338 11943
rect 9366 11690 9394 11695
rect 9310 11689 9394 11690
rect 9310 11663 9367 11689
rect 9393 11663 9394 11689
rect 9310 11662 9394 11663
rect 8862 11657 8890 11662
rect 9366 11657 9394 11662
rect 9254 11634 9282 11639
rect 9254 11633 9338 11634
rect 9254 11607 9255 11633
rect 9281 11607 9338 11633
rect 9254 11606 9338 11607
rect 9254 11601 9282 11606
rect 8750 11578 8778 11583
rect 8750 11531 8778 11550
rect 8918 11577 8946 11583
rect 8918 11551 8919 11577
rect 8945 11551 8946 11577
rect 8918 11410 8946 11551
rect 8918 11377 8946 11382
rect 8974 11578 9002 11583
rect 8750 11354 8778 11359
rect 8750 11186 8778 11326
rect 8918 11186 8946 11191
rect 8750 11153 8778 11158
rect 8806 11185 8946 11186
rect 8806 11159 8919 11185
rect 8945 11159 8946 11185
rect 8806 11158 8946 11159
rect 8974 11186 9002 11550
rect 9030 11577 9058 11583
rect 9030 11551 9031 11577
rect 9057 11551 9058 11577
rect 9030 11522 9058 11551
rect 9030 11489 9058 11494
rect 9198 11577 9226 11583
rect 9198 11551 9199 11577
rect 9225 11551 9226 11577
rect 9198 11298 9226 11551
rect 9142 11186 9170 11191
rect 8974 11158 9058 11186
rect 8750 11074 8778 11079
rect 8750 11027 8778 11046
rect 8694 10985 8722 10990
rect 8750 10794 8778 10799
rect 8806 10794 8834 11158
rect 8918 11153 8946 11158
rect 8974 11073 9002 11079
rect 8974 11047 8975 11073
rect 9001 11047 9002 11073
rect 8974 11018 9002 11047
rect 8974 10985 9002 10990
rect 8862 10850 8890 10855
rect 8862 10849 8946 10850
rect 8862 10823 8863 10849
rect 8889 10823 8946 10849
rect 8862 10822 8946 10823
rect 8862 10817 8890 10822
rect 8778 10766 8834 10794
rect 8750 10747 8778 10766
rect 8582 10150 8834 10178
rect 8078 10033 8106 10038
rect 8694 10066 8722 10071
rect 8694 10019 8722 10038
rect 8134 9954 8162 9959
rect 7910 9927 7911 9953
rect 7937 9927 7938 9953
rect 7910 9730 7938 9927
rect 7910 9697 7938 9702
rect 8022 9926 8134 9954
rect 7406 9585 7434 9590
rect 8022 9617 8050 9926
rect 8134 9907 8162 9926
rect 8750 9953 8778 9959
rect 8750 9927 8751 9953
rect 8777 9927 8778 9953
rect 8022 9591 8023 9617
rect 8049 9591 8050 9617
rect 8022 9585 8050 9591
rect 8078 9786 8106 9791
rect 7238 9561 7322 9562
rect 7238 9535 7239 9561
rect 7265 9535 7322 9561
rect 7238 9534 7322 9535
rect 7238 9529 7266 9534
rect 7070 9366 7210 9394
rect 7182 9338 7210 9366
rect 7182 9291 7210 9310
rect 7014 9226 7042 9231
rect 6846 9225 7042 9226
rect 6846 9199 7015 9225
rect 7041 9199 7042 9225
rect 6846 9198 7042 9199
rect 6790 9087 6791 9113
rect 6817 9087 6818 9113
rect 6790 9081 6818 9087
rect 7014 8889 7042 9198
rect 7014 8863 7015 8889
rect 7041 8863 7042 8889
rect 7014 8857 7042 8863
rect 6510 8409 6538 8414
rect 6902 8833 6930 8839
rect 6902 8807 6903 8833
rect 6929 8807 6930 8833
rect 6902 8498 6930 8807
rect 7294 8834 7322 9534
rect 7350 9529 7378 9534
rect 8078 9561 8106 9758
rect 8750 9730 8778 9927
rect 8470 9702 8778 9730
rect 8470 9618 8498 9702
rect 8806 9674 8834 10150
rect 8862 10009 8890 10015
rect 8862 9983 8863 10009
rect 8889 9983 8890 10009
rect 8862 9954 8890 9983
rect 8862 9921 8890 9926
rect 8750 9673 8834 9674
rect 8750 9647 8807 9673
rect 8833 9647 8834 9673
rect 8750 9646 8834 9647
rect 8414 9617 8498 9618
rect 8414 9591 8471 9617
rect 8497 9591 8498 9617
rect 8414 9590 8498 9591
rect 8078 9535 8079 9561
rect 8105 9535 8106 9561
rect 8078 9529 8106 9535
rect 8302 9562 8330 9567
rect 8302 9515 8330 9534
rect 8190 9506 8218 9511
rect 7294 8787 7322 8806
rect 8134 9505 8218 9506
rect 8134 9479 8191 9505
rect 8217 9479 8218 9505
rect 8134 9478 8218 9479
rect 6902 8385 6930 8470
rect 7462 8498 7490 8503
rect 7462 8451 7490 8470
rect 7630 8497 7658 8503
rect 7630 8471 7631 8497
rect 7657 8471 7658 8497
rect 6902 8359 6903 8385
rect 6929 8359 6930 8385
rect 6902 8353 6930 8359
rect 7126 8442 7154 8447
rect 7126 8385 7154 8414
rect 7126 8359 7127 8385
rect 7153 8359 7154 8385
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 7014 7658 7042 7663
rect 7126 7658 7154 8359
rect 7350 8330 7378 8335
rect 7350 7713 7378 8302
rect 7630 8274 7658 8471
rect 8078 8498 8106 8503
rect 8134 8498 8162 9478
rect 8190 9473 8218 9478
rect 8358 9338 8386 9343
rect 8358 9291 8386 9310
rect 8414 9281 8442 9590
rect 8470 9585 8498 9590
rect 8694 9618 8722 9623
rect 8694 9571 8722 9590
rect 8750 9506 8778 9646
rect 8806 9641 8834 9646
rect 8918 9898 8946 10822
rect 8918 9617 8946 9870
rect 9030 9618 9058 11158
rect 9142 11139 9170 11158
rect 9086 10066 9114 10071
rect 9086 10009 9114 10038
rect 9086 9983 9087 10009
rect 9113 9983 9114 10009
rect 9086 9977 9114 9983
rect 9198 9954 9226 11270
rect 9254 11074 9282 11079
rect 9254 10793 9282 11046
rect 9254 10767 9255 10793
rect 9281 10767 9282 10793
rect 9254 10761 9282 10767
rect 9142 9926 9226 9954
rect 9254 10009 9282 10015
rect 9254 9983 9255 10009
rect 9281 9983 9282 10009
rect 9086 9898 9114 9903
rect 9142 9898 9170 9926
rect 9086 9897 9170 9898
rect 9086 9871 9087 9897
rect 9113 9871 9170 9897
rect 9086 9870 9170 9871
rect 9086 9865 9114 9870
rect 9254 9842 9282 9983
rect 9254 9809 9282 9814
rect 8918 9591 8919 9617
rect 8945 9591 8946 9617
rect 8918 9585 8946 9591
rect 8974 9617 9058 9618
rect 8974 9591 9031 9617
rect 9057 9591 9058 9617
rect 8974 9590 9058 9591
rect 8414 9255 8415 9281
rect 8441 9255 8442 9281
rect 8414 9249 8442 9255
rect 8638 9478 8778 9506
rect 8358 9114 8386 9119
rect 8078 8497 8162 8498
rect 8078 8471 8079 8497
rect 8105 8471 8162 8497
rect 8078 8470 8162 8471
rect 8302 9113 8386 9114
rect 8302 9087 8359 9113
rect 8385 9087 8386 9113
rect 8302 9086 8386 9087
rect 8302 8553 8330 9086
rect 8358 9081 8386 9086
rect 8302 8527 8303 8553
rect 8329 8527 8330 8553
rect 8078 8465 8106 8470
rect 8190 8441 8218 8447
rect 8190 8415 8191 8441
rect 8217 8415 8218 8441
rect 8190 8386 8218 8415
rect 8190 8353 8218 8358
rect 8134 8330 8162 8335
rect 8134 8283 8162 8302
rect 7630 8241 7658 8246
rect 8302 8049 8330 8527
rect 8302 8023 8303 8049
rect 8329 8023 8330 8049
rect 8302 8017 8330 8023
rect 8414 9058 8442 9063
rect 8414 8274 8442 9030
rect 8638 9002 8666 9478
rect 8974 9450 9002 9590
rect 9030 9585 9058 9590
rect 9142 9786 9170 9791
rect 8694 9422 9002 9450
rect 8694 9281 8722 9422
rect 8694 9255 8695 9281
rect 8721 9255 8722 9281
rect 8694 9249 8722 9255
rect 8806 9225 8834 9231
rect 8806 9199 8807 9225
rect 8833 9199 8834 9225
rect 8806 9058 8834 9199
rect 8806 9025 8834 9030
rect 8638 8969 8666 8974
rect 8918 8497 8946 9422
rect 9142 9337 9170 9758
rect 9142 9311 9143 9337
rect 9169 9311 9170 9337
rect 9142 9305 9170 9311
rect 9254 9506 9282 9511
rect 8974 9226 9002 9231
rect 8974 8553 9002 9198
rect 9086 9226 9114 9231
rect 9254 9226 9282 9478
rect 9310 9338 9338 11606
rect 9422 11018 9450 12726
rect 9478 11914 9506 11919
rect 9478 11867 9506 11886
rect 9702 11858 9730 11863
rect 9702 11811 9730 11830
rect 9478 11578 9506 11583
rect 9478 11129 9506 11550
rect 9758 11522 9786 12950
rect 10150 12698 10178 13119
rect 10654 12698 10682 12703
rect 10150 12697 10682 12698
rect 10150 12671 10655 12697
rect 10681 12671 10682 12697
rect 10150 12670 10682 12671
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12306 9842 12311
rect 9814 12259 9842 12278
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10150 11690 10178 12670
rect 10654 12665 10682 12670
rect 10710 12641 10738 18999
rect 12222 19025 12306 19026
rect 12222 18999 12279 19025
rect 12305 18999 12306 19025
rect 12222 18998 12306 18999
rect 11046 18746 11074 18751
rect 11046 18699 11074 18718
rect 11662 14434 11690 14439
rect 11270 14433 11690 14434
rect 11270 14407 11663 14433
rect 11689 14407 11690 14433
rect 11270 14406 11690 14407
rect 11270 13985 11298 14406
rect 11662 14401 11690 14406
rect 12222 14322 12250 18998
rect 12278 18993 12306 18998
rect 12446 18746 12474 20600
rect 12782 20538 12810 20600
rect 12782 20510 12922 20538
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 12446 18713 12474 18718
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 12614 15106 12642 18607
rect 12894 18354 12922 20510
rect 13118 18970 13146 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 13118 18937 13146 18942
rect 13734 18970 13762 18975
rect 13734 18923 13762 18942
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 12894 18321 12922 18326
rect 13398 18354 13426 18359
rect 13398 18307 13426 18326
rect 12894 18242 12922 18247
rect 12334 15078 12642 15106
rect 12670 18241 12922 18242
rect 12670 18215 12895 18241
rect 12921 18215 12922 18241
rect 12670 18214 12922 18215
rect 12222 14321 12306 14322
rect 12222 14295 12223 14321
rect 12249 14295 12306 14321
rect 12222 14294 12306 14295
rect 12222 14289 12250 14294
rect 11270 13959 11271 13985
rect 11297 13959 11298 13985
rect 11270 13953 11298 13959
rect 11606 14265 11634 14271
rect 11606 14239 11607 14265
rect 11633 14239 11634 14265
rect 10878 13930 10906 13935
rect 10766 13902 10878 13930
rect 10766 13593 10794 13902
rect 10878 13883 10906 13902
rect 11438 13930 11466 13935
rect 10766 13567 10767 13593
rect 10793 13567 10794 13593
rect 10766 13561 10794 13567
rect 11438 13537 11466 13902
rect 11438 13511 11439 13537
rect 11465 13511 11466 13537
rect 11438 13454 11466 13511
rect 11606 13454 11634 14239
rect 11662 14210 11690 14215
rect 11662 14209 11746 14210
rect 11662 14183 11663 14209
rect 11689 14183 11746 14209
rect 11662 14182 11746 14183
rect 11662 14177 11690 14182
rect 11438 13426 11522 13454
rect 10822 12642 10850 12647
rect 10710 12615 10711 12641
rect 10737 12615 10738 12641
rect 10710 12306 10738 12615
rect 10710 12273 10738 12278
rect 10766 12641 10850 12642
rect 10766 12615 10823 12641
rect 10849 12615 10850 12641
rect 10766 12614 10850 12615
rect 10654 11970 10682 11975
rect 10766 11970 10794 12614
rect 10822 12609 10850 12614
rect 11270 12361 11298 12367
rect 11270 12335 11271 12361
rect 11297 12335 11298 12361
rect 10878 12305 10906 12311
rect 10878 12279 10879 12305
rect 10905 12279 10906 12305
rect 10878 12025 10906 12279
rect 11270 12306 11298 12335
rect 11494 12306 11522 13426
rect 11550 13426 11634 13454
rect 11662 13874 11690 13879
rect 11550 13257 11578 13426
rect 11550 13231 11551 13257
rect 11577 13231 11578 13257
rect 11550 13225 11578 13231
rect 11662 13257 11690 13846
rect 11718 13538 11746 14182
rect 12278 13874 12306 14294
rect 12334 14265 12362 15078
rect 12334 14239 12335 14265
rect 12361 14239 12362 14265
rect 12334 14233 12362 14239
rect 12670 14042 12698 18214
rect 12894 18209 12922 18214
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 12670 14041 12922 14042
rect 12670 14015 12671 14041
rect 12697 14015 12922 14041
rect 12670 14014 12922 14015
rect 12670 14009 12698 14014
rect 12614 13929 12642 13935
rect 12614 13903 12615 13929
rect 12641 13903 12642 13929
rect 12334 13874 12362 13879
rect 12306 13873 12362 13874
rect 12306 13847 12335 13873
rect 12361 13847 12362 13873
rect 12306 13846 12362 13847
rect 12278 13827 12306 13846
rect 12334 13841 12362 13846
rect 11998 13818 12026 13823
rect 11718 13510 11802 13538
rect 11662 13231 11663 13257
rect 11689 13231 11690 13257
rect 11662 13225 11690 13231
rect 11718 13454 11746 13459
rect 11718 13258 11746 13426
rect 11718 13201 11746 13230
rect 11718 13175 11719 13201
rect 11745 13175 11746 13201
rect 11718 13169 11746 13175
rect 11774 13090 11802 13510
rect 11830 13481 11858 13487
rect 11830 13455 11831 13481
rect 11857 13455 11858 13481
rect 11830 13257 11858 13455
rect 11830 13231 11831 13257
rect 11857 13231 11858 13257
rect 11830 13225 11858 13231
rect 11270 12305 11522 12306
rect 11270 12279 11495 12305
rect 11521 12279 11522 12305
rect 11270 12278 11522 12279
rect 10878 11999 10879 12025
rect 10905 11999 10906 12025
rect 10878 11993 10906 11999
rect 10654 11969 10794 11970
rect 10654 11943 10655 11969
rect 10681 11943 10794 11969
rect 10654 11942 10794 11943
rect 10654 11937 10682 11942
rect 10150 11657 10178 11662
rect 10374 11914 10402 11919
rect 10374 11689 10402 11886
rect 10822 11914 10850 11919
rect 10766 11858 10794 11863
rect 10822 11858 10850 11886
rect 11382 11914 11410 11919
rect 10766 11857 10850 11858
rect 10766 11831 10767 11857
rect 10793 11831 10850 11857
rect 10766 11830 10850 11831
rect 10878 11857 10906 11863
rect 10878 11831 10879 11857
rect 10905 11831 10906 11857
rect 10766 11825 10794 11830
rect 10374 11663 10375 11689
rect 10401 11663 10402 11689
rect 10374 11657 10402 11663
rect 9926 11633 9954 11639
rect 9926 11607 9927 11633
rect 9953 11607 9954 11633
rect 9870 11577 9898 11583
rect 9870 11551 9871 11577
rect 9897 11551 9898 11577
rect 9870 11522 9898 11551
rect 9646 11494 9898 11522
rect 9590 11186 9618 11191
rect 9478 11103 9479 11129
rect 9505 11103 9506 11129
rect 9478 11097 9506 11103
rect 9534 11185 9618 11186
rect 9534 11159 9591 11185
rect 9617 11159 9618 11185
rect 9534 11158 9618 11159
rect 9478 11018 9506 11023
rect 9422 10990 9478 11018
rect 9366 10066 9394 10071
rect 9366 9617 9394 10038
rect 9478 10010 9506 10990
rect 9478 9977 9506 9982
rect 9366 9591 9367 9617
rect 9393 9591 9394 9617
rect 9366 9585 9394 9591
rect 9534 9842 9562 11158
rect 9590 11153 9618 11158
rect 9310 9305 9338 9310
rect 9534 9281 9562 9814
rect 9590 10010 9618 10015
rect 9590 9337 9618 9982
rect 9646 9561 9674 11494
rect 9926 11298 9954 11607
rect 10038 11578 10066 11583
rect 10038 11531 10066 11550
rect 10486 11577 10514 11583
rect 10486 11551 10487 11577
rect 10513 11551 10514 11577
rect 10318 11522 10346 11527
rect 10346 11494 10402 11522
rect 10318 11475 10346 11494
rect 9702 11270 9954 11298
rect 9702 9786 9730 11270
rect 9814 11186 9842 11191
rect 9814 10906 9842 11158
rect 10262 11185 10290 11191
rect 10262 11159 10263 11185
rect 10289 11159 10290 11185
rect 9870 11074 9898 11093
rect 9870 11041 9898 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9814 10878 9898 10906
rect 9814 10402 9842 10407
rect 9814 10355 9842 10374
rect 9870 10290 9898 10878
rect 10206 10570 10234 10575
rect 10038 10458 10066 10463
rect 10038 10411 10066 10430
rect 10206 10401 10234 10542
rect 10206 10375 10207 10401
rect 10233 10375 10234 10401
rect 10206 10369 10234 10375
rect 9982 10290 10010 10295
rect 9814 10289 10010 10290
rect 9814 10263 9983 10289
rect 10009 10263 10010 10289
rect 9814 10262 10010 10263
rect 9758 9954 9786 9959
rect 9814 9954 9842 10262
rect 9982 10257 10010 10262
rect 10094 10289 10122 10295
rect 10094 10263 10095 10289
rect 10121 10263 10122 10289
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10094 10066 10122 10263
rect 10094 10033 10122 10038
rect 10262 10066 10290 11159
rect 10318 11130 10346 11135
rect 10318 11083 10346 11102
rect 9982 10010 10010 10015
rect 10262 10010 10290 10038
rect 10374 10066 10402 11494
rect 10486 11298 10514 11551
rect 10486 11265 10514 11270
rect 10822 10737 10850 10743
rect 10822 10711 10823 10737
rect 10849 10711 10850 10737
rect 10822 10402 10850 10711
rect 10822 10355 10850 10374
rect 10878 10122 10906 11831
rect 10822 10094 10906 10122
rect 10934 11802 10962 11807
rect 10374 10065 10458 10066
rect 10374 10039 10375 10065
rect 10401 10039 10458 10065
rect 10374 10038 10458 10039
rect 10374 10033 10402 10038
rect 9982 9963 10010 9982
rect 10150 10009 10290 10010
rect 10150 9983 10263 10009
rect 10289 9983 10290 10009
rect 10150 9982 10290 9983
rect 9786 9926 9842 9954
rect 9758 9907 9786 9926
rect 9702 9753 9730 9758
rect 9646 9535 9647 9561
rect 9673 9535 9674 9561
rect 9646 9529 9674 9535
rect 9702 9617 9730 9623
rect 9926 9618 9954 9623
rect 9702 9591 9703 9617
rect 9729 9591 9730 9617
rect 9590 9311 9591 9337
rect 9617 9311 9618 9337
rect 9590 9305 9618 9311
rect 9702 9506 9730 9591
rect 9534 9255 9535 9281
rect 9561 9255 9562 9281
rect 9534 9249 9562 9255
rect 9086 9225 9282 9226
rect 9086 9199 9087 9225
rect 9113 9199 9282 9225
rect 9086 9198 9282 9199
rect 9366 9226 9394 9231
rect 9086 9193 9114 9198
rect 9366 9179 9394 9198
rect 9310 9170 9338 9175
rect 9310 9123 9338 9142
rect 9702 8722 9730 9478
rect 9814 9617 9954 9618
rect 9814 9591 9927 9617
rect 9953 9591 9954 9617
rect 9814 9590 9954 9591
rect 9758 9225 9786 9231
rect 9758 9199 9759 9225
rect 9785 9199 9786 9225
rect 9758 9170 9786 9199
rect 9814 9226 9842 9590
rect 9926 9585 9954 9590
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10150 9281 10178 9982
rect 10262 9977 10290 9982
rect 10374 9786 10402 9791
rect 10318 9617 10346 9623
rect 10318 9591 10319 9617
rect 10345 9591 10346 9617
rect 10318 9338 10346 9591
rect 10374 9561 10402 9758
rect 10430 9618 10458 10038
rect 10710 10065 10738 10071
rect 10710 10039 10711 10065
rect 10737 10039 10738 10065
rect 10542 10010 10570 10015
rect 10542 9963 10570 9982
rect 10710 9786 10738 10039
rect 10822 9898 10850 10094
rect 10878 10010 10906 10015
rect 10878 9963 10906 9982
rect 10934 9953 10962 11774
rect 11046 11298 11074 11303
rect 11046 11185 11074 11270
rect 11046 11159 11047 11185
rect 11073 11159 11074 11185
rect 11046 11153 11074 11159
rect 11214 11130 11242 11135
rect 11242 11102 11354 11130
rect 11214 11083 11242 11102
rect 11158 11074 11186 11079
rect 11102 11073 11186 11074
rect 11102 11047 11159 11073
rect 11185 11047 11186 11073
rect 11102 11046 11186 11047
rect 11102 10122 11130 11046
rect 11158 11041 11186 11046
rect 11102 10066 11130 10094
rect 11102 10065 11186 10066
rect 11102 10039 11103 10065
rect 11129 10039 11186 10065
rect 11102 10038 11186 10039
rect 11102 10033 11130 10038
rect 10934 9927 10935 9953
rect 10961 9927 10962 9953
rect 10934 9921 10962 9927
rect 10990 10009 11018 10015
rect 10990 9983 10991 10009
rect 11017 9983 11018 10009
rect 10990 9898 11018 9983
rect 10822 9870 10906 9898
rect 10710 9753 10738 9758
rect 10430 9585 10458 9590
rect 10766 9618 10794 9637
rect 10766 9585 10794 9590
rect 10374 9535 10375 9561
rect 10401 9535 10402 9561
rect 10374 9506 10402 9535
rect 10374 9473 10402 9478
rect 10822 9506 10850 9511
rect 10822 9459 10850 9478
rect 10878 9394 10906 9870
rect 11018 9870 11074 9898
rect 10766 9366 10906 9394
rect 10934 9505 10962 9511
rect 10934 9479 10935 9505
rect 10961 9479 10962 9505
rect 10934 9394 10962 9479
rect 10430 9338 10458 9343
rect 10318 9337 10458 9338
rect 10318 9311 10431 9337
rect 10457 9311 10458 9337
rect 10318 9310 10458 9311
rect 10150 9255 10151 9281
rect 10177 9255 10178 9281
rect 10150 9249 10178 9255
rect 9814 9193 9842 9198
rect 9870 9225 9898 9231
rect 9870 9199 9871 9225
rect 9897 9199 9898 9225
rect 9758 8834 9786 9142
rect 9870 9114 9898 9199
rect 10318 9226 10346 9231
rect 10318 9179 10346 9198
rect 9898 9086 10010 9114
rect 9870 9081 9898 9086
rect 9926 8834 9954 8839
rect 9758 8833 9954 8834
rect 9758 8807 9927 8833
rect 9953 8807 9954 8833
rect 9758 8806 9954 8807
rect 9926 8801 9954 8806
rect 9982 8777 10010 9086
rect 10374 9058 10402 9310
rect 10430 9305 10458 9310
rect 10486 9338 10514 9343
rect 10486 9169 10514 9310
rect 10486 9143 10487 9169
rect 10513 9143 10514 9169
rect 10486 9137 10514 9143
rect 10766 9170 10794 9366
rect 10934 9361 10962 9366
rect 10766 9137 10794 9142
rect 10822 9281 10850 9287
rect 10822 9255 10823 9281
rect 10849 9255 10850 9281
rect 10374 9025 10402 9030
rect 9982 8751 9983 8777
rect 10009 8751 10010 8777
rect 9982 8745 10010 8751
rect 10206 9002 10234 9007
rect 9758 8722 9786 8727
rect 9702 8694 9758 8722
rect 8974 8527 8975 8553
rect 9001 8527 9002 8553
rect 8974 8521 9002 8527
rect 9758 8553 9786 8694
rect 10094 8721 10122 8727
rect 10094 8695 10095 8721
rect 10121 8695 10122 8721
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10094 8610 10122 8695
rect 10094 8577 10122 8582
rect 9758 8527 9759 8553
rect 9785 8527 9786 8553
rect 9758 8521 9786 8527
rect 10150 8554 10178 8559
rect 10150 8507 10178 8526
rect 10206 8553 10234 8974
rect 10766 8778 10794 8783
rect 10766 8731 10794 8750
rect 10206 8527 10207 8553
rect 10233 8527 10234 8553
rect 10206 8521 10234 8527
rect 10598 8721 10626 8727
rect 10598 8695 10599 8721
rect 10625 8695 10626 8721
rect 10598 8554 10626 8695
rect 10710 8722 10738 8727
rect 10710 8675 10738 8694
rect 10822 8610 10850 9255
rect 10878 9282 10906 9287
rect 10990 9282 11018 9870
rect 11046 9729 11074 9870
rect 11046 9703 11047 9729
rect 11073 9703 11074 9729
rect 11046 9697 11074 9703
rect 11158 9561 11186 10038
rect 11270 10009 11298 10015
rect 11270 9983 11271 10009
rect 11297 9983 11298 10009
rect 11270 9954 11298 9983
rect 11270 9921 11298 9926
rect 11214 9674 11242 9679
rect 11214 9673 11298 9674
rect 11214 9647 11215 9673
rect 11241 9647 11298 9673
rect 11214 9646 11298 9647
rect 11214 9641 11242 9646
rect 11158 9535 11159 9561
rect 11185 9535 11186 9561
rect 11158 9529 11186 9535
rect 11270 9506 11298 9646
rect 11158 9394 11186 9399
rect 10878 9281 11018 9282
rect 10878 9255 10879 9281
rect 10905 9255 11018 9281
rect 10878 9254 11018 9255
rect 11046 9282 11074 9287
rect 10878 9249 10906 9254
rect 10878 9170 10906 9175
rect 10878 9113 10906 9142
rect 10878 9087 10879 9113
rect 10905 9087 10906 9113
rect 10878 8722 10906 9087
rect 11046 8945 11074 9254
rect 11046 8919 11047 8945
rect 11073 8919 11074 8945
rect 11046 8913 11074 8919
rect 10878 8689 10906 8694
rect 10990 8833 11018 8839
rect 10990 8807 10991 8833
rect 11017 8807 11018 8833
rect 10822 8577 10850 8582
rect 10598 8521 10626 8526
rect 10990 8554 11018 8807
rect 11046 8722 11074 8727
rect 11046 8675 11074 8694
rect 10990 8521 11018 8526
rect 8918 8471 8919 8497
rect 8945 8471 8946 8497
rect 8918 8465 8946 8471
rect 9590 8497 9618 8503
rect 9590 8471 9591 8497
rect 9617 8471 9618 8497
rect 8694 8442 8722 8447
rect 8414 8049 8442 8246
rect 8414 8023 8415 8049
rect 8441 8023 8442 8049
rect 8414 8017 8442 8023
rect 8470 8441 8722 8442
rect 8470 8415 8695 8441
rect 8721 8415 8722 8441
rect 8470 8414 8722 8415
rect 7350 7687 7351 7713
rect 7377 7687 7378 7713
rect 7350 7681 7378 7687
rect 8358 7937 8386 7943
rect 8358 7911 8359 7937
rect 8385 7911 8386 7937
rect 7014 7657 7154 7658
rect 7014 7631 7015 7657
rect 7041 7631 7154 7657
rect 7014 7630 7154 7631
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7014 7322 7042 7630
rect 8358 7574 8386 7911
rect 8022 7546 8386 7574
rect 8414 7601 8442 7607
rect 8414 7575 8415 7601
rect 8441 7575 8442 7601
rect 8414 7574 8442 7575
rect 8470 7574 8498 8414
rect 8694 8409 8722 8414
rect 9086 8441 9114 8447
rect 9086 8415 9087 8441
rect 9113 8415 9114 8441
rect 8918 8386 8946 8391
rect 8918 8339 8946 8358
rect 8638 8049 8666 8055
rect 8638 8023 8639 8049
rect 8665 8023 8666 8049
rect 8638 7770 8666 8023
rect 8862 7770 8890 7775
rect 8638 7769 8890 7770
rect 8638 7743 8863 7769
rect 8889 7743 8890 7769
rect 8638 7742 8890 7743
rect 8862 7737 8890 7742
rect 9030 7770 9058 7775
rect 9030 7723 9058 7742
rect 8918 7713 8946 7719
rect 8918 7687 8919 7713
rect 8945 7687 8946 7713
rect 8414 7546 8498 7574
rect 8750 7601 8778 7607
rect 8750 7575 8751 7601
rect 8777 7575 8778 7601
rect 7014 7289 7042 7294
rect 7686 7322 7714 7327
rect 7686 7265 7714 7294
rect 8022 7321 8050 7546
rect 8022 7295 8023 7321
rect 8049 7295 8050 7321
rect 8022 7289 8050 7295
rect 7686 7239 7687 7265
rect 7713 7239 7714 7265
rect 7686 7233 7714 7239
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8414 4242 8442 7546
rect 8750 7322 8778 7575
rect 8918 7322 8946 7687
rect 9086 7658 9114 8415
rect 9422 7938 9450 7943
rect 9198 7658 9226 7663
rect 9086 7657 9226 7658
rect 9086 7631 9199 7657
rect 9225 7631 9226 7657
rect 9086 7630 9226 7631
rect 9198 7602 9226 7630
rect 9422 7657 9450 7910
rect 9422 7631 9423 7657
rect 9449 7631 9450 7657
rect 9422 7625 9450 7631
rect 9198 7569 9226 7574
rect 9590 7602 9618 8471
rect 10318 8442 10346 8447
rect 10318 8395 10346 8414
rect 10430 8442 10458 8447
rect 10430 8441 10626 8442
rect 10430 8415 10431 8441
rect 10457 8415 10626 8441
rect 10430 8414 10626 8415
rect 10430 8409 10458 8414
rect 10262 8385 10290 8391
rect 10262 8359 10263 8385
rect 10289 8359 10290 8385
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9758 7714 9786 7719
rect 9758 7667 9786 7686
rect 10262 7714 10290 8359
rect 10598 8049 10626 8414
rect 10598 8023 10599 8049
rect 10625 8023 10626 8049
rect 10598 8017 10626 8023
rect 10710 8078 10850 8106
rect 10710 7993 10738 8078
rect 10710 7967 10711 7993
rect 10737 7967 10738 7993
rect 10710 7961 10738 7967
rect 10766 7993 10794 7999
rect 10766 7967 10767 7993
rect 10793 7967 10794 7993
rect 10262 7681 10290 7686
rect 9590 7569 9618 7574
rect 10766 7602 10794 7967
rect 9086 7322 9114 7327
rect 8918 7321 9114 7322
rect 8918 7295 9087 7321
rect 9113 7295 9114 7321
rect 8918 7294 9114 7295
rect 8750 7289 8778 7294
rect 9086 6426 9114 7294
rect 9310 7322 9338 7327
rect 9310 7275 9338 7294
rect 10766 7266 10794 7574
rect 10710 7238 10794 7266
rect 10822 7601 10850 8078
rect 10990 7938 11018 7943
rect 10990 7891 11018 7910
rect 11158 7714 11186 9366
rect 11158 7667 11186 7686
rect 11270 7713 11298 9478
rect 11326 9337 11354 11102
rect 11382 9730 11410 11886
rect 11494 11858 11522 12278
rect 11718 13062 11802 13090
rect 11942 13201 11970 13207
rect 11942 13175 11943 13201
rect 11969 13175 11970 13201
rect 11662 11970 11690 11975
rect 11662 11923 11690 11942
rect 11494 11825 11522 11830
rect 11550 11913 11578 11919
rect 11550 11887 11551 11913
rect 11577 11887 11578 11913
rect 11550 11690 11578 11887
rect 11718 11858 11746 13062
rect 11942 11970 11970 13175
rect 11998 13201 12026 13790
rect 12614 13482 12642 13903
rect 12670 13818 12698 13823
rect 12670 13771 12698 13790
rect 12894 13593 12922 14014
rect 13006 13930 13034 13935
rect 13034 13902 13146 13930
rect 13006 13883 13034 13902
rect 12894 13567 12895 13593
rect 12921 13567 12922 13593
rect 12894 13561 12922 13567
rect 13118 13593 13146 13902
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13118 13567 13119 13593
rect 13145 13567 13146 13593
rect 13118 13561 13146 13567
rect 12614 13449 12642 13454
rect 11998 13175 11999 13201
rect 12025 13175 12026 13201
rect 11998 13169 12026 13175
rect 13006 13146 13034 13151
rect 12782 12754 12810 12759
rect 12950 12754 12978 12759
rect 12810 12753 12978 12754
rect 12810 12727 12951 12753
rect 12977 12727 12978 12753
rect 12810 12726 12978 12727
rect 12782 12707 12810 12726
rect 12950 12721 12978 12726
rect 13006 12697 13034 13118
rect 13006 12671 13007 12697
rect 13033 12671 13034 12697
rect 13006 12665 13034 12671
rect 13398 13146 13426 13151
rect 12222 12642 12250 12647
rect 12222 12473 12250 12614
rect 12614 12642 12642 12647
rect 12614 12595 12642 12614
rect 12726 12641 12754 12647
rect 12726 12615 12727 12641
rect 12753 12615 12754 12641
rect 12222 12447 12223 12473
rect 12249 12447 12250 12473
rect 12222 12441 12250 12447
rect 12054 12361 12082 12367
rect 12054 12335 12055 12361
rect 12081 12335 12082 12361
rect 11774 11858 11802 11863
rect 11718 11857 11802 11858
rect 11718 11831 11775 11857
rect 11801 11831 11802 11857
rect 11718 11830 11802 11831
rect 11774 11802 11802 11830
rect 11774 11769 11802 11774
rect 11830 11857 11858 11863
rect 11830 11831 11831 11857
rect 11857 11831 11858 11857
rect 11830 11746 11858 11831
rect 11830 11713 11858 11718
rect 11494 11662 11578 11690
rect 11718 11690 11746 11695
rect 11438 11521 11466 11527
rect 11438 11495 11439 11521
rect 11465 11495 11466 11521
rect 11438 11298 11466 11495
rect 11494 11354 11522 11662
rect 11718 11643 11746 11662
rect 11886 11578 11914 11583
rect 11886 11531 11914 11550
rect 11550 11522 11578 11527
rect 11550 11475 11578 11494
rect 11494 11321 11522 11326
rect 11438 11265 11466 11270
rect 11886 10906 11914 10911
rect 11942 10906 11970 11942
rect 11998 11969 12026 11975
rect 11998 11943 11999 11969
rect 12025 11943 12026 11969
rect 11998 11858 12026 11943
rect 12054 11914 12082 12335
rect 12110 12362 12138 12367
rect 12334 12362 12362 12367
rect 12110 12361 12194 12362
rect 12110 12335 12111 12361
rect 12137 12335 12194 12361
rect 12110 12334 12194 12335
rect 12110 12329 12138 12334
rect 12054 11881 12082 11886
rect 12110 12138 12138 12143
rect 11998 11825 12026 11830
rect 11998 11746 12026 11751
rect 11998 11689 12026 11718
rect 11998 11663 11999 11689
rect 12025 11663 12026 11689
rect 11998 11657 12026 11663
rect 12110 11577 12138 12110
rect 12110 11551 12111 11577
rect 12137 11551 12138 11577
rect 12110 11545 12138 11551
rect 12110 11354 12138 11359
rect 12166 11354 12194 12334
rect 12222 12361 12362 12362
rect 12222 12335 12335 12361
rect 12361 12335 12362 12361
rect 12222 12334 12362 12335
rect 12222 11690 12250 12334
rect 12334 12329 12362 12334
rect 12670 12361 12698 12367
rect 12670 12335 12671 12361
rect 12697 12335 12698 12361
rect 12390 12306 12418 12311
rect 12390 12259 12418 12278
rect 12222 11577 12250 11662
rect 12222 11551 12223 11577
rect 12249 11551 12250 11577
rect 12222 11545 12250 11551
rect 12334 11913 12362 11919
rect 12334 11887 12335 11913
rect 12361 11887 12362 11913
rect 12278 11522 12306 11527
rect 12334 11522 12362 11887
rect 12278 11521 12362 11522
rect 12278 11495 12279 11521
rect 12305 11495 12362 11521
rect 12278 11494 12362 11495
rect 12670 11858 12698 12335
rect 12726 12362 12754 12615
rect 12726 12329 12754 12334
rect 13118 12641 13146 12647
rect 13118 12615 13119 12641
rect 13145 12615 13146 12641
rect 13006 12306 13034 12311
rect 13006 12259 13034 12278
rect 13118 12138 13146 12615
rect 13118 12105 13146 12110
rect 13398 12025 13426 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18830 12753 18858 12759
rect 18830 12727 18831 12753
rect 18857 12727 18858 12753
rect 18830 12474 18858 12727
rect 18830 12441 18858 12446
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 14406 12418 14434 12423
rect 14406 12371 14434 12390
rect 14070 12362 14098 12367
rect 14070 12305 14098 12334
rect 14294 12362 14322 12367
rect 14294 12315 14322 12334
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 14070 12279 14071 12305
rect 14097 12279 14098 12305
rect 14070 12273 14098 12279
rect 14630 12305 14658 12311
rect 14630 12279 14631 12305
rect 14657 12279 14658 12305
rect 13398 11999 13399 12025
rect 13425 11999 13426 12025
rect 13398 11993 13426 11999
rect 13622 11970 13650 11975
rect 13622 11923 13650 11942
rect 14630 11970 14658 12279
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 14630 11937 14658 11942
rect 12670 11521 12698 11830
rect 12670 11495 12671 11521
rect 12697 11495 12698 11521
rect 12278 11489 12306 11494
rect 12138 11326 12194 11354
rect 12502 11354 12530 11359
rect 12110 11321 12138 11326
rect 11886 10905 11942 10906
rect 11886 10879 11887 10905
rect 11913 10879 11942 10905
rect 11886 10878 11942 10879
rect 11886 10873 11914 10878
rect 11942 10859 11970 10878
rect 12278 11298 12306 11303
rect 12278 11185 12306 11270
rect 12278 11159 12279 11185
rect 12305 11159 12306 11185
rect 12278 10905 12306 11159
rect 12502 11185 12530 11326
rect 12502 11159 12503 11185
rect 12529 11159 12530 11185
rect 12502 11153 12530 11159
rect 12558 11297 12586 11303
rect 12558 11271 12559 11297
rect 12585 11271 12586 11297
rect 12558 11130 12586 11271
rect 12670 11186 12698 11495
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 14238 11242 14266 11247
rect 12782 11186 12810 11191
rect 12670 11185 12810 11186
rect 12670 11159 12783 11185
rect 12809 11159 12810 11185
rect 12670 11158 12810 11159
rect 12558 11097 12586 11102
rect 12614 11129 12642 11135
rect 12614 11103 12615 11129
rect 12641 11103 12642 11129
rect 12278 10879 12279 10905
rect 12305 10879 12306 10905
rect 12278 10873 12306 10879
rect 12390 11073 12418 11079
rect 12390 11047 12391 11073
rect 12417 11047 12418 11073
rect 12390 10906 12418 11047
rect 12614 10962 12642 11103
rect 12614 10929 12642 10934
rect 12390 10873 12418 10878
rect 12670 10906 12698 10911
rect 12670 10859 12698 10878
rect 11998 10794 12026 10799
rect 12222 10794 12250 10799
rect 11998 10793 12250 10794
rect 11998 10767 11999 10793
rect 12025 10767 12223 10793
rect 12249 10767 12250 10793
rect 11998 10766 12250 10767
rect 11998 10458 12026 10766
rect 12222 10761 12250 10766
rect 12390 10793 12418 10799
rect 12390 10767 12391 10793
rect 12417 10767 12418 10793
rect 11998 10425 12026 10430
rect 11438 10122 11466 10127
rect 11438 10066 11466 10094
rect 11774 10122 11802 10127
rect 11606 10066 11634 10071
rect 11438 10065 11634 10066
rect 11438 10039 11439 10065
rect 11465 10039 11607 10065
rect 11633 10039 11634 10065
rect 11438 10038 11634 10039
rect 11438 10033 11466 10038
rect 11606 10033 11634 10038
rect 11774 10065 11802 10094
rect 11774 10039 11775 10065
rect 11801 10039 11802 10065
rect 11438 9730 11466 9735
rect 11382 9729 11466 9730
rect 11382 9703 11439 9729
rect 11465 9703 11466 9729
rect 11382 9702 11466 9703
rect 11774 9730 11802 10039
rect 12334 10010 12362 10015
rect 12390 10010 12418 10767
rect 12334 10009 12418 10010
rect 12334 9983 12335 10009
rect 12361 9983 12418 10009
rect 12334 9982 12418 9983
rect 12334 9977 12362 9982
rect 12166 9898 12194 9903
rect 12054 9897 12194 9898
rect 12054 9871 12167 9897
rect 12193 9871 12194 9897
rect 12054 9870 12194 9871
rect 11774 9702 11970 9730
rect 11438 9697 11466 9702
rect 11326 9311 11327 9337
rect 11353 9311 11354 9337
rect 11326 9305 11354 9311
rect 11382 9561 11410 9567
rect 11382 9535 11383 9561
rect 11409 9535 11410 9561
rect 11382 8778 11410 9535
rect 11774 9561 11802 9567
rect 11774 9535 11775 9561
rect 11801 9535 11802 9561
rect 11438 9506 11466 9511
rect 11438 9459 11466 9478
rect 11774 9338 11802 9535
rect 11886 9506 11914 9511
rect 11942 9506 11970 9702
rect 12054 9673 12082 9870
rect 12166 9865 12194 9870
rect 12334 9898 12362 9903
rect 12334 9851 12362 9870
rect 12054 9647 12055 9673
rect 12081 9647 12082 9673
rect 12054 9641 12082 9647
rect 11998 9618 12026 9623
rect 11998 9571 12026 9590
rect 12334 9617 12362 9623
rect 12334 9591 12335 9617
rect 12361 9591 12362 9617
rect 12054 9506 12082 9511
rect 11942 9505 12082 9506
rect 11942 9479 12055 9505
rect 12081 9479 12082 9505
rect 11942 9478 12082 9479
rect 11886 9459 11914 9478
rect 11774 9305 11802 9310
rect 11382 8745 11410 8750
rect 11494 9281 11522 9287
rect 11494 9255 11495 9281
rect 11521 9255 11522 9281
rect 11494 8386 11522 9255
rect 11606 8554 11634 8559
rect 11606 8497 11634 8526
rect 11606 8471 11607 8497
rect 11633 8471 11634 8497
rect 11606 8465 11634 8471
rect 11886 8498 11914 8503
rect 11886 8451 11914 8470
rect 11662 8442 11690 8447
rect 11662 8395 11690 8414
rect 11774 8441 11802 8447
rect 11774 8415 11775 8441
rect 11801 8415 11802 8441
rect 11494 8353 11522 8358
rect 11774 8386 11802 8415
rect 11774 8353 11802 8358
rect 11270 7687 11271 7713
rect 11297 7687 11298 7713
rect 11270 7681 11298 7687
rect 11382 7938 11410 7943
rect 10822 7575 10823 7601
rect 10849 7575 10850 7601
rect 10710 7209 10738 7238
rect 10710 7183 10711 7209
rect 10737 7183 10738 7209
rect 10710 7177 10738 7183
rect 10766 7154 10794 7159
rect 10766 7107 10794 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9870 6817 9898 6823
rect 9870 6791 9871 6817
rect 9897 6791 9898 6817
rect 9870 6762 9898 6791
rect 9870 6729 9898 6734
rect 10822 6594 10850 7575
rect 10934 7657 10962 7663
rect 10934 7631 10935 7657
rect 10961 7631 10962 7657
rect 10934 7574 10962 7631
rect 11382 7658 11410 7910
rect 12054 7882 12082 9478
rect 12334 9450 12362 9591
rect 12334 9338 12362 9422
rect 12334 9305 12362 9310
rect 12390 9226 12418 9982
rect 12390 9193 12418 9198
rect 12446 10794 12474 10799
rect 12446 9561 12474 10766
rect 12726 10346 12754 11158
rect 12782 11153 12810 11158
rect 13174 11130 13202 11135
rect 13174 11083 13202 11102
rect 13230 10962 13258 10967
rect 13118 10906 13146 10911
rect 13118 10859 13146 10878
rect 13230 10905 13258 10934
rect 13230 10879 13231 10905
rect 13257 10879 13258 10905
rect 13230 10873 13258 10879
rect 14238 10906 14266 11214
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 14238 10873 14266 10878
rect 12782 10794 12810 10799
rect 12782 10747 12810 10766
rect 12894 10793 12922 10799
rect 12894 10767 12895 10793
rect 12921 10767 12922 10793
rect 12838 10737 12866 10743
rect 12838 10711 12839 10737
rect 12865 10711 12866 10737
rect 12838 10458 12866 10711
rect 12894 10570 12922 10767
rect 12894 10537 12922 10542
rect 13062 10793 13090 10799
rect 13062 10767 13063 10793
rect 13089 10767 13090 10793
rect 12838 10430 12922 10458
rect 12838 10346 12866 10351
rect 12726 10345 12866 10346
rect 12726 10319 12839 10345
rect 12865 10319 12866 10345
rect 12726 10318 12866 10319
rect 12838 10010 12866 10318
rect 12894 10066 12922 10430
rect 13062 10122 13090 10767
rect 20006 10794 20034 11215
rect 20006 10761 20034 10766
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 13062 10089 13090 10094
rect 12894 10033 12922 10038
rect 13846 10066 13874 10071
rect 13846 10019 13874 10038
rect 12782 9954 12810 9959
rect 12782 9907 12810 9926
rect 12446 9535 12447 9561
rect 12473 9535 12474 9561
rect 12334 9170 12362 9175
rect 12334 9123 12362 9142
rect 12446 9114 12474 9535
rect 12838 9617 12866 9982
rect 14182 10010 14210 10015
rect 14182 9963 14210 9982
rect 13230 9898 13258 9903
rect 13230 9673 13258 9870
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 13230 9647 13231 9673
rect 13257 9647 13258 9673
rect 13230 9641 13258 9647
rect 14294 9673 14322 9679
rect 14294 9647 14295 9673
rect 14321 9647 14322 9673
rect 12838 9591 12839 9617
rect 12865 9591 12866 9617
rect 12670 9506 12698 9511
rect 12838 9506 12866 9591
rect 14294 9618 14322 9647
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 14294 9585 14322 9590
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 12670 9505 12866 9506
rect 12670 9479 12671 9505
rect 12697 9479 12866 9505
rect 12670 9478 12866 9479
rect 12614 9282 12642 9287
rect 12614 9235 12642 9254
rect 12166 8554 12194 8559
rect 12166 8049 12194 8526
rect 12446 8498 12474 9086
rect 12278 8386 12306 8391
rect 12278 8162 12306 8358
rect 12278 8050 12306 8134
rect 12166 8023 12167 8049
rect 12193 8023 12194 8049
rect 12166 8017 12194 8023
rect 12222 8049 12306 8050
rect 12222 8023 12279 8049
rect 12305 8023 12306 8049
rect 12222 8022 12306 8023
rect 12054 7849 12082 7854
rect 12166 7770 12194 7775
rect 11886 7769 12194 7770
rect 11886 7743 12167 7769
rect 12193 7743 12194 7769
rect 11886 7742 12194 7743
rect 11046 7601 11074 7607
rect 11046 7575 11047 7601
rect 11073 7575 11074 7601
rect 11046 7574 11074 7575
rect 10878 7546 10962 7574
rect 10990 7546 11074 7574
rect 10878 7265 10906 7546
rect 10878 7239 10879 7265
rect 10905 7239 10906 7265
rect 10878 7233 10906 7239
rect 8806 6398 9114 6426
rect 10654 6566 10850 6594
rect 10878 7154 10906 7159
rect 10878 6762 10906 7126
rect 10934 6930 10962 6935
rect 10990 6930 11018 7546
rect 10934 6929 11018 6930
rect 10934 6903 10935 6929
rect 10961 6903 11018 6929
rect 10934 6902 11018 6903
rect 11382 7266 11410 7630
rect 11662 7714 11690 7719
rect 11662 7657 11690 7686
rect 11886 7713 11914 7742
rect 12166 7737 12194 7742
rect 11886 7687 11887 7713
rect 11913 7687 11914 7713
rect 11886 7681 11914 7687
rect 11662 7631 11663 7657
rect 11689 7631 11690 7657
rect 11662 7625 11690 7631
rect 11998 7658 12026 7663
rect 12222 7658 12250 8022
rect 12278 8017 12306 8022
rect 12390 8050 12418 8055
rect 12390 8003 12418 8022
rect 12446 8049 12474 8470
rect 12446 8023 12447 8049
rect 12473 8023 12474 8049
rect 12446 8017 12474 8023
rect 12670 9170 12698 9478
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 13006 9338 13034 9343
rect 13006 9337 13314 9338
rect 13006 9311 13007 9337
rect 13033 9311 13314 9337
rect 13006 9310 13314 9311
rect 13006 9305 13034 9310
rect 12670 8722 12698 9142
rect 12726 9225 12754 9231
rect 12726 9199 12727 9225
rect 12753 9199 12754 9225
rect 12726 9114 12754 9199
rect 12894 9226 12922 9245
rect 13230 9226 13258 9231
rect 12894 9193 12922 9198
rect 13118 9225 13258 9226
rect 13118 9199 13231 9225
rect 13257 9199 13258 9225
rect 13118 9198 13258 9199
rect 12726 9081 12754 9086
rect 12894 9114 12922 9119
rect 13118 9114 13146 9198
rect 13230 9193 13258 9198
rect 12894 9113 13146 9114
rect 12894 9087 12895 9113
rect 12921 9087 13146 9113
rect 12894 9086 13146 9087
rect 13174 9114 13202 9119
rect 12894 9081 12922 9086
rect 13174 9067 13202 9086
rect 13230 8890 13258 8895
rect 13286 8890 13314 9310
rect 13230 8889 13314 8890
rect 13230 8863 13231 8889
rect 13257 8863 13314 8889
rect 13230 8862 13314 8863
rect 13342 9225 13370 9231
rect 13342 9199 13343 9225
rect 13369 9199 13370 9225
rect 13342 8890 13370 9199
rect 18942 9225 18970 9231
rect 18942 9199 18943 9225
rect 18969 9199 18970 9225
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 13230 8857 13258 8862
rect 13342 8857 13370 8862
rect 14294 8890 14322 8895
rect 14294 8843 14322 8862
rect 14630 8890 14658 8895
rect 12838 8833 12866 8839
rect 12838 8807 12839 8833
rect 12865 8807 12866 8833
rect 12838 8722 12866 8807
rect 14630 8833 14658 8862
rect 14630 8807 14631 8833
rect 14657 8807 14658 8833
rect 14630 8801 14658 8807
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 12670 8721 12866 8722
rect 12670 8695 12671 8721
rect 12697 8695 12866 8721
rect 12670 8694 12866 8695
rect 14742 8722 14770 8727
rect 12558 7938 12586 7943
rect 12558 7891 12586 7910
rect 12334 7770 12362 7775
rect 12278 7714 12306 7719
rect 12278 7667 12306 7686
rect 12334 7713 12362 7742
rect 12334 7687 12335 7713
rect 12361 7687 12362 7713
rect 12334 7681 12362 7687
rect 11998 7657 12250 7658
rect 11998 7631 11999 7657
rect 12025 7631 12250 7657
rect 11998 7630 12250 7631
rect 12614 7658 12642 7663
rect 12670 7658 12698 8694
rect 14742 8675 14770 8694
rect 18942 8722 18970 9199
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 18942 8689 18970 8694
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 12726 8162 12754 8167
rect 12726 8115 12754 8134
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 12782 8050 12810 8055
rect 12782 8003 12810 8022
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 12838 7937 12866 7943
rect 12838 7911 12839 7937
rect 12865 7911 12866 7937
rect 12642 7630 12698 7658
rect 12782 7714 12810 7719
rect 11998 7625 12026 7630
rect 12614 7611 12642 7630
rect 11774 7601 11802 7607
rect 11774 7575 11775 7601
rect 11801 7575 11802 7601
rect 11774 7546 11802 7575
rect 11718 7518 11802 7546
rect 11718 7321 11746 7518
rect 11718 7295 11719 7321
rect 11745 7295 11746 7321
rect 11718 7289 11746 7295
rect 12782 7321 12810 7686
rect 12838 7602 12866 7911
rect 13006 7938 13034 7943
rect 13006 7713 13034 7910
rect 14294 7770 14322 7775
rect 14294 7723 14322 7742
rect 13006 7687 13007 7713
rect 13033 7687 13034 7713
rect 13006 7681 13034 7687
rect 12838 7569 12866 7574
rect 12950 7658 12978 7663
rect 12782 7295 12783 7321
rect 12809 7295 12810 7321
rect 11382 7265 11578 7266
rect 11382 7239 11383 7265
rect 11409 7239 11578 7265
rect 11382 7238 11578 7239
rect 10934 6897 10962 6902
rect 11326 6874 11354 6879
rect 11382 6874 11410 7238
rect 11550 6985 11578 7238
rect 11550 6959 11551 6985
rect 11577 6959 11578 6985
rect 11550 6953 11578 6959
rect 11326 6873 11410 6874
rect 11326 6847 11327 6873
rect 11353 6847 11410 6873
rect 11326 6846 11410 6847
rect 11326 6841 11354 6846
rect 8526 4242 8554 4247
rect 8414 4214 8526 4242
rect 8526 4209 8554 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8750 2058 8778 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8750 400 8778 2030
rect 8806 1777 8834 6398
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 8862 4242 8890 4247
rect 10654 4214 10682 6566
rect 10878 4214 10906 6734
rect 12782 4214 12810 7295
rect 12950 7322 12978 7630
rect 14070 7658 14098 7663
rect 14070 7601 14098 7630
rect 18830 7658 18858 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18830 7625 18858 7630
rect 14070 7575 14071 7601
rect 14097 7575 14098 7601
rect 14070 7569 14098 7575
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13006 7322 13034 7327
rect 12950 7321 13034 7322
rect 12950 7295 13007 7321
rect 13033 7295 13034 7321
rect 12950 7294 13034 7295
rect 13006 7289 13034 7294
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 8862 2169 8890 4214
rect 10542 4186 10682 4214
rect 10710 4186 10906 4214
rect 12614 4186 12810 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 8862 2143 8863 2169
rect 8889 2143 8890 2169
rect 8862 2137 8890 2143
rect 10542 2169 10570 4186
rect 10542 2143 10543 2169
rect 10569 2143 10570 2169
rect 10542 2137 10570 2143
rect 9366 2058 9394 2063
rect 9366 2011 9394 2030
rect 10430 2058 10458 2063
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 2030
rect 10710 1777 10738 4186
rect 11046 2058 11074 2063
rect 11046 2011 11074 2030
rect 10710 1751 10711 1777
rect 10737 1751 10738 1777
rect 10710 1745 10738 1751
rect 12446 1834 12474 1839
rect 11214 1666 11242 1671
rect 11102 1665 11242 1666
rect 11102 1639 11215 1665
rect 11241 1639 11242 1665
rect 11102 1638 11242 1639
rect 11102 400 11130 1638
rect 11214 1633 11242 1638
rect 12446 400 12474 1806
rect 12614 1777 12642 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 13062 1834 13090 1839
rect 13062 1787 13090 1806
rect 12614 1751 12615 1777
rect 12641 1751 12642 1777
rect 12614 1745 12642 1751
rect 17262 1666 17290 1671
rect 17150 1665 17290 1666
rect 17150 1639 17263 1665
rect 17289 1639 17290 1665
rect 17150 1638 17290 1639
rect 17150 400 17178 1638
rect 17262 1633 17290 1638
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 10416 0 10472 400
rect 11088 0 11144 400
rect 12432 0 12488 400
rect 17136 0 17192 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8750 18718 8778 18746
rect 9366 18745 9394 18746
rect 9366 18719 9367 18745
rect 9367 18719 9393 18745
rect 9393 18719 9394 18745
rect 9366 18718 9394 18719
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2086 13790 2114 13818
rect 966 12446 994 12474
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 11774 994 11802
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 8358 13537 8386 13538
rect 8358 13511 8359 13537
rect 8359 13511 8385 13537
rect 8385 13511 8386 13537
rect 8358 13510 8386 13511
rect 7014 13062 7042 13090
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 4998 12809 5026 12810
rect 4998 12783 4999 12809
rect 4999 12783 5025 12809
rect 5025 12783 5026 12809
rect 4998 12782 5026 12783
rect 6902 12782 6930 12810
rect 2142 12753 2170 12754
rect 2142 12727 2143 12753
rect 2143 12727 2169 12753
rect 2169 12727 2170 12753
rect 2142 12726 2170 12727
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 5502 12305 5530 12306
rect 5502 12279 5503 12305
rect 5503 12279 5529 12305
rect 5529 12279 5530 12305
rect 5502 12278 5530 12279
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 5502 12054 5530 12082
rect 6454 12614 6482 12642
rect 6790 12054 6818 12082
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 6454 11969 6482 11970
rect 6454 11943 6455 11969
rect 6455 11943 6481 11969
rect 6481 11943 6482 11969
rect 6454 11942 6482 11943
rect 9590 14406 9618 14434
rect 9310 14182 9338 14210
rect 9254 13929 9282 13930
rect 9254 13903 9255 13929
rect 9255 13903 9281 13929
rect 9281 13903 9282 13929
rect 9254 13902 9282 13903
rect 8526 13537 8554 13538
rect 8526 13511 8527 13537
rect 8527 13511 8553 13537
rect 8553 13511 8554 13537
rect 8526 13510 8554 13511
rect 8582 13062 8610 13090
rect 8638 12753 8666 12754
rect 8638 12727 8639 12753
rect 8639 12727 8665 12753
rect 8665 12727 8666 12753
rect 8638 12726 8666 12727
rect 7350 12670 7378 12698
rect 7966 12697 7994 12698
rect 7966 12671 7967 12697
rect 7967 12671 7993 12697
rect 7993 12671 7994 12697
rect 7966 12670 7994 12671
rect 7014 12641 7042 12642
rect 7014 12615 7015 12641
rect 7015 12615 7041 12641
rect 7041 12615 7042 12641
rect 7014 12614 7042 12615
rect 8134 12446 8162 12474
rect 8694 12473 8722 12474
rect 8694 12447 8695 12473
rect 8695 12447 8721 12473
rect 8721 12447 8722 12473
rect 8694 12446 8722 12447
rect 6902 11942 6930 11970
rect 6902 11774 6930 11802
rect 7574 12025 7602 12026
rect 7574 11999 7575 12025
rect 7575 11999 7601 12025
rect 7601 11999 7602 12025
rect 7574 11998 7602 11999
rect 6846 11577 6874 11578
rect 6846 11551 6847 11577
rect 6847 11551 6873 11577
rect 6873 11551 6874 11577
rect 6846 11550 6874 11551
rect 7014 11494 7042 11522
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6734 11382 6762 11410
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 4998 11158 5026 11186
rect 2086 11046 2114 11074
rect 966 10766 994 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 7014 11382 7042 11410
rect 6902 11129 6930 11130
rect 6902 11103 6903 11129
rect 6903 11103 6929 11129
rect 6929 11103 6930 11129
rect 6902 11102 6930 11103
rect 6062 10934 6090 10962
rect 6790 10934 6818 10962
rect 6454 10430 6482 10458
rect 4998 10374 5026 10402
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 5334 9673 5362 9674
rect 5334 9647 5335 9673
rect 5335 9647 5361 9673
rect 5361 9647 5362 9673
rect 5334 9646 5362 9647
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 6398 9590 6426 9618
rect 6062 9198 6090 9226
rect 6006 9169 6034 9170
rect 6006 9143 6007 9169
rect 6007 9143 6033 9169
rect 6033 9143 6034 9169
rect 6006 9142 6034 9143
rect 6454 9142 6482 9170
rect 6286 9086 6314 9114
rect 6454 8470 6482 8498
rect 4998 8414 5026 8442
rect 5502 8441 5530 8442
rect 5502 8415 5503 8441
rect 5503 8415 5529 8441
rect 5529 8415 5530 8441
rect 5502 8414 5530 8415
rect 6790 10457 6818 10458
rect 6790 10431 6791 10457
rect 6791 10431 6817 10457
rect 6817 10431 6818 10457
rect 6790 10430 6818 10431
rect 6734 10374 6762 10402
rect 6846 10038 6874 10066
rect 6678 9926 6706 9954
rect 7182 11494 7210 11522
rect 7182 11214 7210 11242
rect 7070 10065 7098 10066
rect 7070 10039 7071 10065
rect 7071 10039 7097 10065
rect 7097 10039 7098 10065
rect 7070 10038 7098 10039
rect 7126 11102 7154 11130
rect 7014 10009 7042 10010
rect 7014 9983 7015 10009
rect 7015 9983 7041 10009
rect 7041 9983 7042 10009
rect 7014 9982 7042 9983
rect 7350 11185 7378 11186
rect 7350 11159 7351 11185
rect 7351 11159 7377 11185
rect 7377 11159 7378 11185
rect 7350 11158 7378 11159
rect 7406 10766 7434 10794
rect 7798 10934 7826 10962
rect 7294 10430 7322 10458
rect 6902 9870 6930 9898
rect 7014 9729 7042 9730
rect 7014 9703 7015 9729
rect 7015 9703 7041 9729
rect 7041 9703 7042 9729
rect 7014 9702 7042 9703
rect 6566 9225 6594 9226
rect 6566 9199 6567 9225
rect 6567 9199 6593 9225
rect 6593 9199 6594 9225
rect 6566 9198 6594 9199
rect 6734 9086 6762 9114
rect 6846 9617 6874 9618
rect 6846 9591 6847 9617
rect 6847 9591 6873 9617
rect 6873 9591 6874 9617
rect 6846 9590 6874 9591
rect 7350 9982 7378 10010
rect 7294 9953 7322 9954
rect 7294 9927 7295 9953
rect 7295 9927 7321 9953
rect 7321 9927 7322 9953
rect 7294 9926 7322 9927
rect 7182 9673 7210 9674
rect 7182 9647 7183 9673
rect 7183 9647 7209 9673
rect 7209 9647 7210 9673
rect 7182 9646 7210 9647
rect 7406 10038 7434 10066
rect 7910 10542 7938 10570
rect 7462 9953 7490 9954
rect 7462 9927 7463 9953
rect 7463 9927 7489 9953
rect 7489 9927 7490 9953
rect 7462 9926 7490 9927
rect 7966 10457 7994 10458
rect 7966 10431 7967 10457
rect 7967 10431 7993 10457
rect 7993 10431 7994 10457
rect 7966 10430 7994 10431
rect 8190 10934 8218 10962
rect 8414 10793 8442 10794
rect 8414 10767 8415 10793
rect 8415 10767 8441 10793
rect 8441 10767 8442 10793
rect 8414 10766 8442 10767
rect 8806 11998 8834 12026
rect 8638 11913 8666 11914
rect 8638 11887 8639 11913
rect 8639 11887 8665 11913
rect 8665 11887 8666 11913
rect 8638 11886 8666 11887
rect 8694 11718 8722 11746
rect 9030 11830 9058 11858
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 12110 19110 12138 19138
rect 10430 18718 10458 18746
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9926 14433 9954 14434
rect 9926 14407 9927 14433
rect 9927 14407 9953 14433
rect 9953 14407 9954 14433
rect 9926 14406 9954 14407
rect 9814 14294 9842 14322
rect 10094 14209 10122 14210
rect 10094 14183 10095 14209
rect 10095 14183 10121 14209
rect 10121 14183 10122 14209
rect 10094 14182 10122 14183
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9982 14014 10010 14042
rect 10206 14265 10234 14266
rect 10206 14239 10207 14265
rect 10207 14239 10233 14265
rect 10233 14239 10234 14265
rect 10206 14238 10234 14239
rect 10206 14014 10234 14042
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 10318 13257 10346 13258
rect 10318 13231 10319 13257
rect 10319 13231 10345 13257
rect 10345 13231 10346 13257
rect 10318 13230 10346 13231
rect 9422 12726 9450 12754
rect 9198 11942 9226 11970
rect 9254 11913 9282 11914
rect 9254 11887 9255 11913
rect 9255 11887 9281 11913
rect 9281 11887 9282 11913
rect 9254 11886 9282 11887
rect 8750 11577 8778 11578
rect 8750 11551 8751 11577
rect 8751 11551 8777 11577
rect 8777 11551 8778 11577
rect 8750 11550 8778 11551
rect 8918 11382 8946 11410
rect 8974 11550 9002 11578
rect 8750 11326 8778 11354
rect 8750 11158 8778 11186
rect 9030 11494 9058 11522
rect 9198 11270 9226 11298
rect 8750 11073 8778 11074
rect 8750 11047 8751 11073
rect 8751 11047 8777 11073
rect 8777 11047 8778 11073
rect 8750 11046 8778 11047
rect 8694 10990 8722 11018
rect 8974 10990 9002 11018
rect 8750 10793 8778 10794
rect 8750 10767 8751 10793
rect 8751 10767 8777 10793
rect 8777 10767 8778 10793
rect 8750 10766 8778 10767
rect 8078 10038 8106 10066
rect 8694 10065 8722 10066
rect 8694 10039 8695 10065
rect 8695 10039 8721 10065
rect 8721 10039 8722 10065
rect 8694 10038 8722 10039
rect 7910 9702 7938 9730
rect 8134 9953 8162 9954
rect 8134 9927 8135 9953
rect 8135 9927 8161 9953
rect 8161 9927 8162 9953
rect 8134 9926 8162 9927
rect 7406 9590 7434 9618
rect 8078 9758 8106 9786
rect 7182 9337 7210 9338
rect 7182 9311 7183 9337
rect 7183 9311 7209 9337
rect 7209 9311 7210 9337
rect 7182 9310 7210 9311
rect 6510 8414 6538 8442
rect 7350 9534 7378 9562
rect 8862 9926 8890 9954
rect 8302 9561 8330 9562
rect 8302 9535 8303 9561
rect 8303 9535 8329 9561
rect 8329 9535 8330 9561
rect 8302 9534 8330 9535
rect 7294 8833 7322 8834
rect 7294 8807 7295 8833
rect 7295 8807 7321 8833
rect 7321 8807 7322 8833
rect 7294 8806 7322 8807
rect 6902 8470 6930 8498
rect 7462 8497 7490 8498
rect 7462 8471 7463 8497
rect 7463 8471 7489 8497
rect 7489 8471 7490 8497
rect 7462 8470 7490 8471
rect 7126 8414 7154 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 7350 8302 7378 8330
rect 8358 9337 8386 9338
rect 8358 9311 8359 9337
rect 8359 9311 8385 9337
rect 8385 9311 8386 9337
rect 8358 9310 8386 9311
rect 8694 9617 8722 9618
rect 8694 9591 8695 9617
rect 8695 9591 8721 9617
rect 8721 9591 8722 9617
rect 8694 9590 8722 9591
rect 8918 9870 8946 9898
rect 9142 11185 9170 11186
rect 9142 11159 9143 11185
rect 9143 11159 9169 11185
rect 9169 11159 9170 11185
rect 9142 11158 9170 11159
rect 9086 10038 9114 10066
rect 9254 11046 9282 11074
rect 9254 9814 9282 9842
rect 8190 8358 8218 8386
rect 8134 8329 8162 8330
rect 8134 8303 8135 8329
rect 8135 8303 8161 8329
rect 8161 8303 8162 8329
rect 8134 8302 8162 8303
rect 7630 8246 7658 8274
rect 8414 9030 8442 9058
rect 9142 9758 9170 9786
rect 8806 9030 8834 9058
rect 8638 8974 8666 9002
rect 9254 9505 9282 9506
rect 9254 9479 9255 9505
rect 9255 9479 9281 9505
rect 9281 9479 9282 9505
rect 9254 9478 9282 9479
rect 8974 9225 9002 9226
rect 8974 9199 8975 9225
rect 8975 9199 9001 9225
rect 9001 9199 9002 9225
rect 8974 9198 9002 9199
rect 9478 11913 9506 11914
rect 9478 11887 9479 11913
rect 9479 11887 9505 11913
rect 9505 11887 9506 11913
rect 9478 11886 9506 11887
rect 9702 11857 9730 11858
rect 9702 11831 9703 11857
rect 9703 11831 9729 11857
rect 9729 11831 9730 11857
rect 9702 11830 9730 11831
rect 9478 11550 9506 11578
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9814 12305 9842 12306
rect 9814 12279 9815 12305
rect 9815 12279 9841 12305
rect 9841 12279 9842 12305
rect 9814 12278 9842 12279
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 11046 18745 11074 18746
rect 11046 18719 11047 18745
rect 11047 18719 11073 18745
rect 11073 18719 11074 18745
rect 11046 18718 11074 18719
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 12446 18718 12474 18746
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 13118 18942 13146 18970
rect 13734 18969 13762 18970
rect 13734 18943 13735 18969
rect 13735 18943 13761 18969
rect 13761 18943 13762 18969
rect 13734 18942 13762 18943
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 12894 18326 12922 18354
rect 13398 18353 13426 18354
rect 13398 18327 13399 18353
rect 13399 18327 13425 18353
rect 13425 18327 13426 18353
rect 13398 18326 13426 18327
rect 10878 13929 10906 13930
rect 10878 13903 10879 13929
rect 10879 13903 10905 13929
rect 10905 13903 10906 13929
rect 10878 13902 10906 13903
rect 11438 13902 11466 13930
rect 10710 12278 10738 12306
rect 11662 13846 11690 13874
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 12278 13846 12306 13874
rect 11998 13790 12026 13818
rect 11718 13426 11746 13454
rect 11718 13230 11746 13258
rect 10150 11662 10178 11690
rect 10374 11886 10402 11914
rect 10822 11886 10850 11914
rect 11382 11886 11410 11914
rect 9478 10990 9506 11018
rect 9366 10038 9394 10066
rect 9478 9982 9506 10010
rect 9534 9814 9562 9842
rect 9310 9310 9338 9338
rect 9590 9982 9618 10010
rect 10038 11577 10066 11578
rect 10038 11551 10039 11577
rect 10039 11551 10065 11577
rect 10065 11551 10066 11577
rect 10038 11550 10066 11551
rect 10318 11521 10346 11522
rect 10318 11495 10319 11521
rect 10319 11495 10345 11521
rect 10345 11495 10346 11521
rect 10318 11494 10346 11495
rect 9814 11185 9842 11186
rect 9814 11159 9815 11185
rect 9815 11159 9841 11185
rect 9841 11159 9842 11185
rect 9814 11158 9842 11159
rect 9870 11073 9898 11074
rect 9870 11047 9871 11073
rect 9871 11047 9897 11073
rect 9897 11047 9898 11073
rect 9870 11046 9898 11047
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9814 10401 9842 10402
rect 9814 10375 9815 10401
rect 9815 10375 9841 10401
rect 9841 10375 9842 10401
rect 9814 10374 9842 10375
rect 10206 10542 10234 10570
rect 10038 10457 10066 10458
rect 10038 10431 10039 10457
rect 10039 10431 10065 10457
rect 10065 10431 10066 10457
rect 10038 10430 10066 10431
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10094 10038 10122 10066
rect 10318 11129 10346 11130
rect 10318 11103 10319 11129
rect 10319 11103 10345 11129
rect 10345 11103 10346 11129
rect 10318 11102 10346 11103
rect 10262 10038 10290 10066
rect 10486 11270 10514 11298
rect 10822 10401 10850 10402
rect 10822 10375 10823 10401
rect 10823 10375 10849 10401
rect 10849 10375 10850 10401
rect 10822 10374 10850 10375
rect 10934 11774 10962 11802
rect 9982 10009 10010 10010
rect 9982 9983 9983 10009
rect 9983 9983 10009 10009
rect 10009 9983 10010 10009
rect 9982 9982 10010 9983
rect 9758 9953 9786 9954
rect 9758 9927 9759 9953
rect 9759 9927 9785 9953
rect 9785 9927 9786 9953
rect 9758 9926 9786 9927
rect 9702 9758 9730 9786
rect 9702 9478 9730 9506
rect 9366 9225 9394 9226
rect 9366 9199 9367 9225
rect 9367 9199 9393 9225
rect 9393 9199 9394 9225
rect 9366 9198 9394 9199
rect 9310 9169 9338 9170
rect 9310 9143 9311 9169
rect 9311 9143 9337 9169
rect 9337 9143 9338 9169
rect 9310 9142 9338 9143
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10374 9758 10402 9786
rect 10542 10009 10570 10010
rect 10542 9983 10543 10009
rect 10543 9983 10569 10009
rect 10569 9983 10570 10009
rect 10542 9982 10570 9983
rect 10878 10009 10906 10010
rect 10878 9983 10879 10009
rect 10879 9983 10905 10009
rect 10905 9983 10906 10009
rect 10878 9982 10906 9983
rect 11046 11270 11074 11298
rect 11214 11129 11242 11130
rect 11214 11103 11215 11129
rect 11215 11103 11241 11129
rect 11241 11103 11242 11129
rect 11214 11102 11242 11103
rect 11102 10094 11130 10122
rect 10710 9758 10738 9786
rect 10430 9590 10458 9618
rect 10766 9617 10794 9618
rect 10766 9591 10767 9617
rect 10767 9591 10793 9617
rect 10793 9591 10794 9617
rect 10766 9590 10794 9591
rect 10374 9478 10402 9506
rect 10822 9505 10850 9506
rect 10822 9479 10823 9505
rect 10823 9479 10849 9505
rect 10849 9479 10850 9505
rect 10822 9478 10850 9479
rect 10990 9870 11018 9898
rect 10934 9366 10962 9394
rect 9814 9198 9842 9226
rect 9758 9142 9786 9170
rect 10318 9225 10346 9226
rect 10318 9199 10319 9225
rect 10319 9199 10345 9225
rect 10345 9199 10346 9225
rect 10318 9198 10346 9199
rect 9870 9086 9898 9114
rect 10486 9310 10514 9338
rect 10766 9142 10794 9170
rect 10374 9030 10402 9058
rect 10206 8974 10234 9002
rect 9758 8694 9786 8722
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10094 8582 10122 8610
rect 10150 8553 10178 8554
rect 10150 8527 10151 8553
rect 10151 8527 10177 8553
rect 10177 8527 10178 8553
rect 10150 8526 10178 8527
rect 10766 8777 10794 8778
rect 10766 8751 10767 8777
rect 10767 8751 10793 8777
rect 10793 8751 10794 8777
rect 10766 8750 10794 8751
rect 10710 8721 10738 8722
rect 10710 8695 10711 8721
rect 10711 8695 10737 8721
rect 10737 8695 10738 8721
rect 10710 8694 10738 8695
rect 11270 9926 11298 9954
rect 11270 9478 11298 9506
rect 11158 9366 11186 9394
rect 11046 9254 11074 9282
rect 10878 9142 10906 9170
rect 10878 8694 10906 8722
rect 10822 8582 10850 8610
rect 10598 8526 10626 8554
rect 11046 8721 11074 8722
rect 11046 8695 11047 8721
rect 11047 8695 11073 8721
rect 11073 8695 11074 8721
rect 11046 8694 11074 8695
rect 10990 8526 11018 8554
rect 8414 8246 8442 8274
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8918 8385 8946 8386
rect 8918 8359 8919 8385
rect 8919 8359 8945 8385
rect 8945 8359 8946 8385
rect 8918 8358 8946 8359
rect 9030 7769 9058 7770
rect 9030 7743 9031 7769
rect 9031 7743 9057 7769
rect 9057 7743 9058 7769
rect 9030 7742 9058 7743
rect 7014 7294 7042 7322
rect 7686 7294 7714 7322
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 8750 7294 8778 7322
rect 9422 7910 9450 7938
rect 9198 7574 9226 7602
rect 10318 8441 10346 8442
rect 10318 8415 10319 8441
rect 10319 8415 10345 8441
rect 10345 8415 10346 8441
rect 10318 8414 10346 8415
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9758 7713 9786 7714
rect 9758 7687 9759 7713
rect 9759 7687 9785 7713
rect 9785 7687 9786 7713
rect 9758 7686 9786 7687
rect 10262 7686 10290 7714
rect 9590 7574 9618 7602
rect 10766 7574 10794 7602
rect 9310 7321 9338 7322
rect 9310 7295 9311 7321
rect 9311 7295 9337 7321
rect 9337 7295 9338 7321
rect 9310 7294 9338 7295
rect 10990 7937 11018 7938
rect 10990 7911 10991 7937
rect 10991 7911 11017 7937
rect 11017 7911 11018 7937
rect 10990 7910 11018 7911
rect 11158 7713 11186 7714
rect 11158 7687 11159 7713
rect 11159 7687 11185 7713
rect 11185 7687 11186 7713
rect 11158 7686 11186 7687
rect 11662 11969 11690 11970
rect 11662 11943 11663 11969
rect 11663 11943 11689 11969
rect 11689 11943 11690 11969
rect 11662 11942 11690 11943
rect 11494 11830 11522 11858
rect 12670 13817 12698 13818
rect 12670 13791 12671 13817
rect 12671 13791 12697 13817
rect 12697 13791 12698 13817
rect 12670 13790 12698 13791
rect 13006 13929 13034 13930
rect 13006 13903 13007 13929
rect 13007 13903 13033 13929
rect 13033 13903 13034 13929
rect 13006 13902 13034 13903
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12614 13454 12642 13482
rect 13006 13118 13034 13146
rect 12782 12753 12810 12754
rect 12782 12727 12783 12753
rect 12783 12727 12809 12753
rect 12809 12727 12810 12753
rect 12782 12726 12810 12727
rect 13398 13118 13426 13146
rect 12222 12614 12250 12642
rect 12614 12641 12642 12642
rect 12614 12615 12615 12641
rect 12615 12615 12641 12641
rect 12641 12615 12642 12641
rect 12614 12614 12642 12615
rect 11942 11942 11970 11970
rect 11774 11774 11802 11802
rect 11830 11718 11858 11746
rect 11718 11689 11746 11690
rect 11718 11663 11719 11689
rect 11719 11663 11745 11689
rect 11745 11663 11746 11689
rect 11718 11662 11746 11663
rect 11886 11577 11914 11578
rect 11886 11551 11887 11577
rect 11887 11551 11913 11577
rect 11913 11551 11914 11577
rect 11886 11550 11914 11551
rect 11550 11521 11578 11522
rect 11550 11495 11551 11521
rect 11551 11495 11577 11521
rect 11577 11495 11578 11521
rect 11550 11494 11578 11495
rect 11494 11326 11522 11354
rect 11438 11270 11466 11298
rect 12054 11886 12082 11914
rect 12110 12110 12138 12138
rect 11998 11830 12026 11858
rect 11998 11718 12026 11746
rect 12390 12305 12418 12306
rect 12390 12279 12391 12305
rect 12391 12279 12417 12305
rect 12417 12279 12418 12305
rect 12390 12278 12418 12279
rect 12222 11662 12250 11690
rect 12726 12334 12754 12362
rect 13006 12305 13034 12306
rect 13006 12279 13007 12305
rect 13007 12279 13033 12305
rect 13033 12279 13034 12305
rect 13006 12278 13034 12279
rect 13118 12110 13146 12138
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 19950 12782 19978 12810
rect 18830 12446 18858 12474
rect 20006 12446 20034 12474
rect 14406 12417 14434 12418
rect 14406 12391 14407 12417
rect 14407 12391 14433 12417
rect 14433 12391 14434 12417
rect 14406 12390 14434 12391
rect 14070 12334 14098 12362
rect 14294 12361 14322 12362
rect 14294 12335 14295 12361
rect 14295 12335 14321 12361
rect 14321 12335 14322 12361
rect 14294 12334 14322 12335
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 13622 11969 13650 11970
rect 13622 11943 13623 11969
rect 13623 11943 13649 11969
rect 13649 11943 13650 11969
rect 13622 11942 13650 11943
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 14630 11942 14658 11970
rect 12670 11830 12698 11858
rect 12110 11326 12138 11354
rect 12502 11326 12530 11354
rect 11942 10878 11970 10906
rect 12278 11270 12306 11298
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14238 11241 14266 11242
rect 14238 11215 14239 11241
rect 14239 11215 14265 11241
rect 14265 11215 14266 11241
rect 14238 11214 14266 11215
rect 12558 11102 12586 11130
rect 12614 10934 12642 10962
rect 12390 10878 12418 10906
rect 12670 10905 12698 10906
rect 12670 10879 12671 10905
rect 12671 10879 12697 10905
rect 12697 10879 12698 10905
rect 12670 10878 12698 10879
rect 11998 10430 12026 10458
rect 11438 10094 11466 10122
rect 11774 10094 11802 10122
rect 11438 9505 11466 9506
rect 11438 9479 11439 9505
rect 11439 9479 11465 9505
rect 11465 9479 11466 9505
rect 11438 9478 11466 9479
rect 11886 9505 11914 9506
rect 11886 9479 11887 9505
rect 11887 9479 11913 9505
rect 11913 9479 11914 9505
rect 11886 9478 11914 9479
rect 12334 9897 12362 9898
rect 12334 9871 12335 9897
rect 12335 9871 12361 9897
rect 12361 9871 12362 9897
rect 12334 9870 12362 9871
rect 11998 9617 12026 9618
rect 11998 9591 11999 9617
rect 11999 9591 12025 9617
rect 12025 9591 12026 9617
rect 11998 9590 12026 9591
rect 11774 9310 11802 9338
rect 11382 8750 11410 8778
rect 11606 8526 11634 8554
rect 11886 8497 11914 8498
rect 11886 8471 11887 8497
rect 11887 8471 11913 8497
rect 11913 8471 11914 8497
rect 11886 8470 11914 8471
rect 11662 8441 11690 8442
rect 11662 8415 11663 8441
rect 11663 8415 11689 8441
rect 11689 8415 11690 8441
rect 11662 8414 11690 8415
rect 11494 8358 11522 8386
rect 11774 8358 11802 8386
rect 11382 7910 11410 7938
rect 10766 7153 10794 7154
rect 10766 7127 10767 7153
rect 10767 7127 10793 7153
rect 10793 7127 10794 7153
rect 10766 7126 10794 7127
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9870 6734 9898 6762
rect 12334 9422 12362 9450
rect 12334 9310 12362 9338
rect 12390 9198 12418 9226
rect 12446 10766 12474 10794
rect 13174 11129 13202 11130
rect 13174 11103 13175 11129
rect 13175 11103 13201 11129
rect 13201 11103 13202 11129
rect 13174 11102 13202 11103
rect 13230 10934 13258 10962
rect 13118 10905 13146 10906
rect 13118 10879 13119 10905
rect 13119 10879 13145 10905
rect 13145 10879 13146 10905
rect 13118 10878 13146 10879
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 14238 10878 14266 10906
rect 12782 10793 12810 10794
rect 12782 10767 12783 10793
rect 12783 10767 12809 10793
rect 12809 10767 12810 10793
rect 12782 10766 12810 10767
rect 12894 10542 12922 10570
rect 20006 10766 20034 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 13062 10094 13090 10122
rect 12894 10038 12922 10066
rect 13846 10065 13874 10066
rect 13846 10039 13847 10065
rect 13847 10039 13873 10065
rect 13873 10039 13874 10065
rect 13846 10038 13874 10039
rect 12838 9982 12866 10010
rect 12782 9953 12810 9954
rect 12782 9927 12783 9953
rect 12783 9927 12809 9953
rect 12809 9927 12810 9953
rect 12782 9926 12810 9927
rect 12334 9169 12362 9170
rect 12334 9143 12335 9169
rect 12335 9143 12361 9169
rect 12361 9143 12362 9169
rect 12334 9142 12362 9143
rect 14182 10009 14210 10010
rect 14182 9983 14183 10009
rect 14183 9983 14209 10009
rect 14209 9983 14210 10009
rect 14182 9982 14210 9983
rect 13230 9870 13258 9898
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14294 9590 14322 9618
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 12614 9281 12642 9282
rect 12614 9255 12615 9281
rect 12615 9255 12641 9281
rect 12641 9255 12642 9281
rect 12614 9254 12642 9255
rect 12446 9086 12474 9114
rect 12166 8526 12194 8554
rect 12446 8470 12474 8498
rect 12278 8358 12306 8386
rect 12278 8134 12306 8162
rect 12054 7854 12082 7882
rect 11382 7630 11410 7658
rect 10878 7126 10906 7154
rect 11662 7686 11690 7714
rect 12390 8049 12418 8050
rect 12390 8023 12391 8049
rect 12391 8023 12417 8049
rect 12417 8023 12418 8049
rect 12390 8022 12418 8023
rect 20006 9422 20034 9450
rect 12670 9142 12698 9170
rect 12894 9225 12922 9226
rect 12894 9199 12895 9225
rect 12895 9199 12921 9225
rect 12921 9199 12922 9225
rect 12894 9198 12922 9199
rect 12726 9086 12754 9114
rect 13174 9113 13202 9114
rect 13174 9087 13175 9113
rect 13175 9087 13201 9113
rect 13201 9087 13202 9113
rect 13174 9086 13202 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 13342 8862 13370 8890
rect 14294 8889 14322 8890
rect 14294 8863 14295 8889
rect 14295 8863 14321 8889
rect 14321 8863 14322 8889
rect 14294 8862 14322 8863
rect 14630 8862 14658 8890
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 14742 8721 14770 8722
rect 14742 8695 14743 8721
rect 14743 8695 14769 8721
rect 14769 8695 14770 8721
rect 14742 8694 14770 8695
rect 12558 7937 12586 7938
rect 12558 7911 12559 7937
rect 12559 7911 12585 7937
rect 12585 7911 12586 7937
rect 12558 7910 12586 7911
rect 12334 7742 12362 7770
rect 12278 7713 12306 7714
rect 12278 7687 12279 7713
rect 12279 7687 12305 7713
rect 12305 7687 12306 7713
rect 12278 7686 12306 7687
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 20006 8750 20034 8778
rect 18942 8694 18970 8722
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 12726 8161 12754 8162
rect 12726 8135 12727 8161
rect 12727 8135 12753 8161
rect 12753 8135 12754 8161
rect 12726 8134 12754 8135
rect 12782 8049 12810 8050
rect 12782 8023 12783 8049
rect 12783 8023 12809 8049
rect 12809 8023 12810 8049
rect 12782 8022 12810 8023
rect 12614 7657 12642 7658
rect 12614 7631 12615 7657
rect 12615 7631 12641 7657
rect 12641 7631 12642 7657
rect 12614 7630 12642 7631
rect 12782 7686 12810 7714
rect 13006 7910 13034 7938
rect 14294 7769 14322 7770
rect 14294 7743 14295 7769
rect 14295 7743 14321 7769
rect 14321 7743 14322 7769
rect 14294 7742 14322 7743
rect 12838 7574 12866 7602
rect 12950 7630 12978 7658
rect 10878 6734 10906 6762
rect 8526 4214 8554 4242
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8750 2030 8778 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 8862 4214 8890 4242
rect 14070 7630 14098 7658
rect 20006 7742 20034 7770
rect 18830 7630 18858 7658
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9366 2057 9394 2058
rect 9366 2031 9367 2057
rect 9367 2031 9393 2057
rect 9393 2031 9394 2057
rect 9366 2030 9394 2031
rect 10430 2030 10458 2058
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11046 2057 11074 2058
rect 11046 2031 11047 2057
rect 11047 2031 11073 2057
rect 11073 2031 11074 2057
rect 11046 2030 11074 2031
rect 12446 1806 12474 1834
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 13062 1833 13090 1834
rect 13062 1807 13063 1833
rect 13063 1807 13089 1833
rect 13089 1807 13090 1833
rect 13062 1806 13090 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 13113 18942 13118 18970
rect 13146 18942 13734 18970
rect 13762 18942 13767 18970
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8745 18718 8750 18746
rect 8778 18718 9366 18746
rect 9394 18718 9399 18746
rect 10425 18718 10430 18746
rect 10458 18718 11046 18746
rect 11074 18718 11079 18746
rect 12441 18718 12446 18746
rect 12474 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 12889 18326 12894 18354
rect 12922 18326 13398 18354
rect 13426 18326 13431 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9585 14406 9590 14434
rect 9618 14406 9926 14434
rect 9954 14406 9959 14434
rect 9809 14294 9814 14322
rect 9842 14294 9847 14322
rect 9814 14266 9842 14294
rect 9814 14238 10206 14266
rect 10234 14238 10239 14266
rect 9305 14182 9310 14210
rect 9338 14182 10094 14210
rect 10122 14182 10127 14210
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 9977 14014 9982 14042
rect 10010 14014 10206 14042
rect 10234 14014 10239 14042
rect 9249 13902 9254 13930
rect 9282 13902 10878 13930
rect 10906 13902 11438 13930
rect 11466 13902 13006 13930
rect 13034 13902 13039 13930
rect 11657 13846 11662 13874
rect 11690 13846 12278 13874
rect 12306 13846 12311 13874
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 11993 13790 11998 13818
rect 12026 13790 12670 13818
rect 12698 13790 12703 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 8353 13510 8358 13538
rect 8386 13510 8526 13538
rect 8554 13510 8559 13538
rect 11718 13454 12614 13482
rect 12642 13454 12647 13482
rect 11713 13426 11718 13454
rect 11746 13426 11751 13454
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 10313 13230 10318 13258
rect 10346 13230 11718 13258
rect 11746 13230 11751 13258
rect 13001 13118 13006 13146
rect 13034 13118 13398 13146
rect 13426 13118 18830 13146
rect 18858 13118 18863 13146
rect 7009 13062 7014 13090
rect 7042 13062 8582 13090
rect 8610 13062 8615 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 20600 12810 21000 12824
rect 4186 12782 4998 12810
rect 5026 12782 6902 12810
rect 6930 12782 6935 12810
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 4186 12754 4214 12782
rect 20600 12768 21000 12782
rect 2137 12726 2142 12754
rect 2170 12726 4214 12754
rect 8633 12726 8638 12754
rect 8666 12726 9422 12754
rect 9450 12726 12782 12754
rect 12810 12726 12815 12754
rect 7345 12670 7350 12698
rect 7378 12670 7966 12698
rect 7994 12670 7999 12698
rect 6449 12614 6454 12642
rect 6482 12614 7014 12642
rect 7042 12614 7047 12642
rect 12217 12614 12222 12642
rect 12250 12614 12614 12642
rect 12642 12614 12647 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 20600 12474 21000 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 8129 12446 8134 12474
rect 8162 12446 8694 12474
rect 8722 12446 8727 12474
rect 15946 12446 18830 12474
rect 18858 12446 18863 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 0 12432 400 12446
rect 15946 12418 15974 12446
rect 20600 12432 21000 12446
rect 14401 12390 14406 12418
rect 14434 12390 15974 12418
rect 2137 12334 2142 12362
rect 2170 12334 4214 12362
rect 12721 12334 12726 12362
rect 12754 12334 14070 12362
rect 14098 12334 14294 12362
rect 14322 12334 18830 12362
rect 18858 12334 18863 12362
rect 4186 12306 4214 12334
rect 4186 12278 5502 12306
rect 5530 12278 5535 12306
rect 9809 12278 9814 12306
rect 9842 12278 10710 12306
rect 10738 12278 10743 12306
rect 12385 12278 12390 12306
rect 12418 12278 13006 12306
rect 13034 12278 13039 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 0 12110 994 12138
rect 12105 12110 12110 12138
rect 12138 12110 13118 12138
rect 13146 12110 13151 12138
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 0 12096 400 12110
rect 20600 12096 21000 12110
rect 5497 12054 5502 12082
rect 5530 12054 6790 12082
rect 6818 12054 6823 12082
rect 4186 11998 7574 12026
rect 7602 11998 8806 12026
rect 8834 11998 8839 12026
rect 4186 11970 4214 11998
rect 2137 11942 2142 11970
rect 2170 11942 4214 11970
rect 6449 11942 6454 11970
rect 6482 11942 6902 11970
rect 6930 11942 6935 11970
rect 9193 11942 9198 11970
rect 9226 11942 9506 11970
rect 11657 11942 11662 11970
rect 11690 11942 11942 11970
rect 11970 11942 11975 11970
rect 13426 11942 13622 11970
rect 13650 11942 14630 11970
rect 14658 11942 14663 11970
rect 9478 11914 9506 11942
rect 8633 11886 8638 11914
rect 8666 11886 9254 11914
rect 9282 11886 9287 11914
rect 9473 11886 9478 11914
rect 9506 11886 10374 11914
rect 10402 11886 10407 11914
rect 10817 11886 10822 11914
rect 10850 11886 11382 11914
rect 11410 11886 12054 11914
rect 12082 11886 12087 11914
rect 13426 11858 13454 11942
rect 9025 11830 9030 11858
rect 9058 11830 9702 11858
rect 9730 11830 11494 11858
rect 11522 11830 11998 11858
rect 12026 11830 12670 11858
rect 12698 11830 13454 11858
rect 0 11802 400 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 6897 11774 6902 11802
rect 6930 11774 6935 11802
rect 10929 11774 10934 11802
rect 10962 11774 11774 11802
rect 11802 11774 11807 11802
rect 0 11760 400 11774
rect 6902 11746 6930 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 6902 11718 8694 11746
rect 8722 11718 8727 11746
rect 11825 11718 11830 11746
rect 11858 11718 11998 11746
rect 12026 11718 12031 11746
rect 6902 11578 6930 11718
rect 8694 11690 8722 11718
rect 8694 11662 10150 11690
rect 10178 11662 10183 11690
rect 11713 11662 11718 11690
rect 11746 11662 12222 11690
rect 12250 11662 12255 11690
rect 6841 11550 6846 11578
rect 6874 11550 6930 11578
rect 8745 11550 8750 11578
rect 8778 11550 8974 11578
rect 9002 11550 9478 11578
rect 9506 11550 9511 11578
rect 10033 11550 10038 11578
rect 10066 11550 11886 11578
rect 11914 11550 11919 11578
rect 7009 11494 7014 11522
rect 7042 11494 7182 11522
rect 7210 11494 7215 11522
rect 9025 11494 9030 11522
rect 9058 11494 10318 11522
rect 10346 11494 11550 11522
rect 11578 11494 11583 11522
rect 6729 11382 6734 11410
rect 6762 11382 7014 11410
rect 7042 11382 8918 11410
rect 8946 11382 8951 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 8745 11326 8750 11354
rect 8778 11326 11494 11354
rect 11522 11326 12110 11354
rect 12138 11326 12502 11354
rect 12530 11326 12535 11354
rect 7546 11270 9198 11298
rect 9226 11270 9231 11298
rect 10481 11270 10486 11298
rect 10514 11270 11046 11298
rect 11074 11270 11438 11298
rect 11466 11270 12278 11298
rect 12306 11270 12311 11298
rect 7546 11242 7574 11270
rect 7177 11214 7182 11242
rect 7210 11214 7574 11242
rect 14233 11214 14238 11242
rect 14266 11214 15974 11242
rect 15946 11186 15974 11214
rect 2137 11158 2142 11186
rect 2170 11158 4998 11186
rect 5026 11158 5031 11186
rect 7345 11158 7350 11186
rect 7378 11158 8750 11186
rect 8778 11158 8783 11186
rect 9137 11158 9142 11186
rect 9170 11158 9814 11186
rect 9842 11158 9847 11186
rect 15946 11158 18830 11186
rect 18858 11158 18863 11186
rect 6897 11102 6902 11130
rect 6930 11102 7126 11130
rect 7154 11102 7159 11130
rect 9366 11102 10318 11130
rect 10346 11102 11214 11130
rect 11242 11102 11247 11130
rect 12553 11102 12558 11130
rect 12586 11102 13174 11130
rect 13202 11102 13207 11130
rect 2081 11046 2086 11074
rect 2114 11046 8750 11074
rect 8778 11046 9254 11074
rect 9282 11046 9287 11074
rect 8689 10990 8694 11018
rect 8722 10990 8974 11018
rect 9002 10990 9007 11018
rect 9366 10962 9394 11102
rect 9478 11046 9870 11074
rect 9898 11046 9903 11074
rect 9478 11018 9506 11046
rect 9473 10990 9478 11018
rect 9506 10990 9511 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 6057 10934 6062 10962
rect 6090 10934 6790 10962
rect 6818 10934 6823 10962
rect 7793 10934 7798 10962
rect 7826 10934 8190 10962
rect 8218 10934 9394 10962
rect 12609 10934 12614 10962
rect 12642 10934 13230 10962
rect 13258 10934 13263 10962
rect 11937 10878 11942 10906
rect 11970 10878 12390 10906
rect 12418 10878 12670 10906
rect 12698 10878 12703 10906
rect 13113 10878 13118 10906
rect 13146 10878 14238 10906
rect 14266 10878 14271 10906
rect 0 10794 400 10808
rect 20600 10794 21000 10808
rect 0 10766 966 10794
rect 994 10766 999 10794
rect 7401 10766 7406 10794
rect 7434 10766 7938 10794
rect 8409 10766 8414 10794
rect 8442 10766 8750 10794
rect 8778 10766 8783 10794
rect 12441 10766 12446 10794
rect 12474 10766 12782 10794
rect 12810 10766 12815 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 0 10752 400 10766
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 7910 10570 7938 10766
rect 20600 10752 21000 10766
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7905 10542 7910 10570
rect 7938 10542 10206 10570
rect 10234 10542 12894 10570
rect 12922 10542 12927 10570
rect 6449 10430 6454 10458
rect 6482 10430 6790 10458
rect 6818 10430 7294 10458
rect 7322 10430 7966 10458
rect 7994 10430 7999 10458
rect 10033 10430 10038 10458
rect 10066 10430 11998 10458
rect 12026 10430 12031 10458
rect 4993 10374 4998 10402
rect 5026 10374 6734 10402
rect 6762 10374 6767 10402
rect 9809 10374 9814 10402
rect 9842 10374 10822 10402
rect 10850 10374 10855 10402
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 11097 10094 11102 10122
rect 11130 10094 11438 10122
rect 11466 10094 11471 10122
rect 11769 10094 11774 10122
rect 11802 10094 13062 10122
rect 13090 10094 13095 10122
rect 6841 10038 6846 10066
rect 6874 10038 7070 10066
rect 7098 10038 7406 10066
rect 7434 10038 7439 10066
rect 8073 10038 8078 10066
rect 8106 10038 8694 10066
rect 8722 10038 9086 10066
rect 9114 10038 9366 10066
rect 9394 10038 10094 10066
rect 10122 10038 10127 10066
rect 10257 10038 10262 10066
rect 10290 10038 10906 10066
rect 12889 10038 12894 10066
rect 12922 10038 13846 10066
rect 13874 10038 13879 10066
rect 10878 10010 10906 10038
rect 7009 9982 7014 10010
rect 7042 9982 7350 10010
rect 7378 9982 7383 10010
rect 8750 9982 9478 10010
rect 9506 9982 9511 10010
rect 9585 9982 9590 10010
rect 9618 9982 9982 10010
rect 10010 9982 10542 10010
rect 10570 9982 10575 10010
rect 10873 9982 10878 10010
rect 10906 9982 10911 10010
rect 12833 9982 12838 10010
rect 12866 9982 14182 10010
rect 14210 9982 14215 10010
rect 6673 9926 6678 9954
rect 6706 9926 7294 9954
rect 7322 9926 7327 9954
rect 7457 9926 7462 9954
rect 7490 9926 8134 9954
rect 8162 9926 8167 9954
rect 8750 9898 8778 9982
rect 8857 9926 8862 9954
rect 8890 9926 9758 9954
rect 9786 9926 9791 9954
rect 11265 9926 11270 9954
rect 11298 9926 12782 9954
rect 12810 9926 12815 9954
rect 6897 9870 6902 9898
rect 6930 9870 8778 9898
rect 8913 9870 8918 9898
rect 8946 9870 10990 9898
rect 11018 9870 11023 9898
rect 11270 9842 11298 9926
rect 12329 9870 12334 9898
rect 12362 9870 13230 9898
rect 13258 9870 13263 9898
rect 9249 9814 9254 9842
rect 9282 9814 9534 9842
rect 9562 9814 11298 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 8073 9758 8078 9786
rect 8106 9758 9142 9786
rect 9170 9758 9702 9786
rect 9730 9758 9735 9786
rect 10369 9758 10374 9786
rect 10402 9758 10710 9786
rect 10738 9758 10743 9786
rect 7009 9702 7014 9730
rect 7042 9702 7910 9730
rect 7938 9702 7943 9730
rect 5329 9646 5334 9674
rect 5362 9646 7182 9674
rect 7210 9646 7215 9674
rect 6393 9590 6398 9618
rect 6426 9590 6846 9618
rect 6874 9590 6879 9618
rect 7401 9590 7406 9618
rect 7434 9590 8694 9618
rect 8722 9590 8727 9618
rect 10425 9590 10430 9618
rect 10458 9590 10766 9618
rect 10794 9590 10799 9618
rect 11993 9590 11998 9618
rect 12026 9590 14294 9618
rect 14322 9590 18830 9618
rect 18858 9590 18863 9618
rect 7345 9534 7350 9562
rect 7378 9534 8302 9562
rect 8330 9534 8335 9562
rect 9249 9478 9254 9506
rect 9282 9478 9702 9506
rect 9730 9478 9735 9506
rect 10369 9478 10374 9506
rect 10402 9478 10822 9506
rect 10850 9478 10855 9506
rect 11265 9478 11270 9506
rect 11298 9478 11438 9506
rect 11466 9478 11886 9506
rect 11914 9478 11919 9506
rect 10822 9450 10850 9478
rect 20600 9450 21000 9464
rect 10822 9422 12334 9450
rect 12362 9422 12367 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 10929 9366 10934 9394
rect 10962 9366 11158 9394
rect 11186 9366 11191 9394
rect 7177 9310 7182 9338
rect 7210 9310 8358 9338
rect 8386 9310 8391 9338
rect 9305 9310 9310 9338
rect 9338 9310 10486 9338
rect 10514 9310 11774 9338
rect 11802 9310 11807 9338
rect 12329 9310 12334 9338
rect 12362 9310 13202 9338
rect 8358 9226 8386 9310
rect 11041 9254 11046 9282
rect 11074 9254 12614 9282
rect 12642 9254 12647 9282
rect 6057 9198 6062 9226
rect 6090 9198 6566 9226
rect 6594 9198 6599 9226
rect 8358 9198 8974 9226
rect 9002 9198 9007 9226
rect 9361 9198 9366 9226
rect 9394 9198 9814 9226
rect 9842 9198 10318 9226
rect 10346 9198 10351 9226
rect 12385 9198 12390 9226
rect 12418 9198 12894 9226
rect 12922 9198 12927 9226
rect 6001 9142 6006 9170
rect 6034 9142 6454 9170
rect 6482 9142 9310 9170
rect 9338 9142 9758 9170
rect 9786 9142 9791 9170
rect 10761 9142 10766 9170
rect 10794 9142 10878 9170
rect 10906 9142 10911 9170
rect 12329 9142 12334 9170
rect 12362 9142 12670 9170
rect 12698 9142 12703 9170
rect 13174 9114 13202 9310
rect 20600 9114 21000 9128
rect 6281 9086 6286 9114
rect 6314 9086 6734 9114
rect 6762 9086 9870 9114
rect 9898 9086 9903 9114
rect 12441 9086 12446 9114
rect 12474 9086 12726 9114
rect 12754 9086 12759 9114
rect 13169 9086 13174 9114
rect 13202 9086 13207 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 8409 9030 8414 9058
rect 8442 9030 8806 9058
rect 8834 9030 10374 9058
rect 10402 9030 10407 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 8633 8974 8638 9002
rect 8666 8974 10206 9002
rect 10234 8974 10239 9002
rect 13337 8862 13342 8890
rect 13370 8862 14294 8890
rect 14322 8862 14630 8890
rect 14658 8862 15974 8890
rect 15946 8834 15974 8862
rect 7289 8806 7294 8834
rect 7322 8806 7574 8834
rect 15946 8806 18830 8834
rect 18858 8806 18863 8834
rect 7546 8778 7574 8806
rect 20600 8778 21000 8792
rect 7546 8750 10766 8778
rect 10794 8750 11382 8778
rect 11410 8750 11415 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 9753 8694 9758 8722
rect 9786 8694 10710 8722
rect 10738 8694 10743 8722
rect 10873 8694 10878 8722
rect 10906 8694 11046 8722
rect 11074 8694 11079 8722
rect 14737 8694 14742 8722
rect 14770 8694 18942 8722
rect 18970 8694 18975 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 10089 8582 10094 8610
rect 10122 8582 10822 8610
rect 10850 8582 11634 8610
rect 11606 8554 11634 8582
rect 10145 8526 10150 8554
rect 10178 8526 10598 8554
rect 10626 8526 10990 8554
rect 11018 8526 11023 8554
rect 11601 8526 11606 8554
rect 11634 8526 12166 8554
rect 12194 8526 12199 8554
rect 6449 8470 6454 8498
rect 6482 8470 6902 8498
rect 6930 8470 7462 8498
rect 7490 8470 7495 8498
rect 11881 8470 11886 8498
rect 11914 8470 12446 8498
rect 12474 8470 12479 8498
rect 4993 8414 4998 8442
rect 5026 8414 5502 8442
rect 5530 8414 6510 8442
rect 6538 8414 7126 8442
rect 7154 8414 7159 8442
rect 10313 8414 10318 8442
rect 10346 8414 11662 8442
rect 11690 8414 11695 8442
rect 8185 8358 8190 8386
rect 8218 8358 8918 8386
rect 8946 8358 8951 8386
rect 11489 8358 11494 8386
rect 11522 8358 11774 8386
rect 11802 8358 12278 8386
rect 12306 8358 12311 8386
rect 7345 8302 7350 8330
rect 7378 8302 8134 8330
rect 8162 8302 8167 8330
rect 7625 8246 7630 8274
rect 7658 8246 8414 8274
rect 8442 8246 8447 8274
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 12273 8134 12278 8162
rect 12306 8134 12726 8162
rect 12754 8134 12759 8162
rect 12385 8022 12390 8050
rect 12418 8022 12782 8050
rect 12810 8022 12815 8050
rect 9417 7910 9422 7938
rect 9450 7910 10990 7938
rect 11018 7910 11382 7938
rect 11410 7910 11415 7938
rect 12553 7910 12558 7938
rect 12586 7910 13006 7938
rect 13034 7910 13039 7938
rect 12049 7854 12054 7882
rect 12082 7854 12087 7882
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 12054 7770 12082 7854
rect 20600 7770 21000 7784
rect 9025 7742 9030 7770
rect 9058 7742 12334 7770
rect 12362 7742 12367 7770
rect 12950 7742 14294 7770
rect 14322 7742 14327 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 9753 7686 9758 7714
rect 9786 7686 10262 7714
rect 10290 7686 10295 7714
rect 11153 7686 11158 7714
rect 11186 7686 11662 7714
rect 11690 7686 11695 7714
rect 12273 7686 12278 7714
rect 12306 7686 12782 7714
rect 12810 7686 12815 7714
rect 12950 7658 12978 7742
rect 20600 7728 21000 7742
rect 11377 7630 11382 7658
rect 11410 7630 12614 7658
rect 12642 7630 12950 7658
rect 12978 7630 12983 7658
rect 13426 7630 14070 7658
rect 14098 7630 18830 7658
rect 18858 7630 18863 7658
rect 13426 7602 13454 7630
rect 9193 7574 9198 7602
rect 9226 7574 9590 7602
rect 9618 7574 10766 7602
rect 10794 7574 10799 7602
rect 12833 7574 12838 7602
rect 12866 7574 13454 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 7009 7294 7014 7322
rect 7042 7294 7686 7322
rect 7714 7294 8750 7322
rect 8778 7294 9310 7322
rect 9338 7294 9343 7322
rect 10761 7126 10766 7154
rect 10794 7126 10878 7154
rect 10906 7126 10911 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 9865 6734 9870 6762
rect 9898 6734 10878 6762
rect 10906 6734 10911 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 8521 4214 8526 4242
rect 8554 4214 8862 4242
rect 8890 4214 8895 4242
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8745 2030 8750 2058
rect 8778 2030 9366 2058
rect 9394 2030 9399 2058
rect 10425 2030 10430 2058
rect 10458 2030 11046 2058
rect 11074 2030 11079 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 12441 1806 12446 1834
rect 12474 1806 13062 1834
rect 13090 1806 13095 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6944 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9464 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10136 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform 1 0 7840 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform -1 0 8568 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform -1 0 6552 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _110_
timestamp 1698175906
transform -1 0 6216 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _111_
timestamp 1698175906
transform -1 0 6384 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6384 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _113_
timestamp 1698175906
transform 1 0 8176 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _114_
timestamp 1698175906
transform -1 0 8512 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _115_
timestamp 1698175906
transform 1 0 9688 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6720 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10304 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform -1 0 12152 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _122_
timestamp 1698175906
transform 1 0 8848 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform 1 0 10080 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform -1 0 12096 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11200 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform -1 0 11312 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform 1 0 12152 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform 1 0 11536 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_
timestamp 1698175906
transform 1 0 10976 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 7392 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1698175906
transform 1 0 9240 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1698175906
transform 1 0 10248 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _135_
timestamp 1698175906
transform 1 0 11704 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform 1 0 12096 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _138_
timestamp 1698175906
transform -1 0 7336 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7560 0 -1 10192
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform -1 0 7560 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform 1 0 10472 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1698175906
transform 1 0 12208 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12992 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 9520 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 10416 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform -1 0 10080 0 1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 12432 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _149_
timestamp 1698175906
transform 1 0 10136 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform 1 0 10696 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform 1 0 11256 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _152_
timestamp 1698175906
transform 1 0 11648 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _153_
timestamp 1698175906
transform -1 0 9520 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _154_
timestamp 1698175906
transform -1 0 7280 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _155_
timestamp 1698175906
transform -1 0 6552 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform 1 0 9128 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698175906
transform -1 0 10360 0 1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 9408 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _159_
timestamp 1698175906
transform -1 0 7224 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _160_
timestamp 1698175906
transform -1 0 6888 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform -1 0 9856 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform 1 0 10640 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _163_
timestamp 1698175906
transform 1 0 10920 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform -1 0 8512 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform -1 0 9744 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9184 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform 1 0 7952 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _169_
timestamp 1698175906
transform 1 0 8008 0 -1 8624
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _170_
timestamp 1698175906
transform -1 0 9128 0 -1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _171_
timestamp 1698175906
transform 1 0 10248 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _172_
timestamp 1698175906
transform 1 0 9128 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _173_
timestamp 1698175906
transform 1 0 10808 0 -1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform -1 0 11816 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698175906
transform 1 0 11536 0 1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _176_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11368 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 12880 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform 1 0 7112 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1698175906
transform 1 0 11312 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11928 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _181_
timestamp 1698175906
transform 1 0 11480 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1698175906
transform 1 0 9800 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform 1 0 12880 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _184_
timestamp 1698175906
transform 1 0 11816 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _185_
timestamp 1698175906
transform 1 0 8456 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _186_
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _187_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9240 0 -1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _188_
timestamp 1698175906
transform -1 0 8232 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform 1 0 9856 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform 1 0 10752 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _191_
timestamp 1698175906
transform -1 0 10864 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform 1 0 10920 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1698175906
transform 1 0 13104 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _194_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _195_
timestamp 1698175906
transform 1 0 12992 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _196_
timestamp 1698175906
transform -1 0 12712 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _197_
timestamp 1698175906
transform -1 0 9240 0 -1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _198_
timestamp 1698175906
transform 1 0 8232 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _199_
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _200_
timestamp 1698175906
transform 1 0 12096 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _202_
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _203_
timestamp 1698175906
transform 1 0 11536 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _204_
timestamp 1698175906
transform -1 0 10864 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _205_
timestamp 1698175906
transform -1 0 10528 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 11368 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 12768 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 5376 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 4872 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 6216 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform -1 0 14336 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 9128 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 11256 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform -1 0 6552 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 8456 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform -1 0 7056 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 11424 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 6888 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform -1 0 9128 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 10808 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 11872 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 6888 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 12768 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 12712 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform -1 0 11368 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 9296 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _233_
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _234_
timestamp 1698175906
transform 1 0 14168 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _235_
timestamp 1698175906
transform 1 0 12096 0 1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6776 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 13104 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 7112 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 7952 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 10752 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 12992 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 7000 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 8344 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 7168 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 11536 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 9688 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform -1 0 13048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 14616 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 13608 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 12656 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 9296 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 11480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 10976 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 8736 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 9912 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 10752 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12432 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 13944 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_290
timestamp 1698175906
transform 1 0 16912 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_294
timestamp 1698175906
transform 1 0 17136 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_299
timestamp 1698175906
transform 1 0 17416 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698175906
transform 1 0 17640 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698175906
transform 1 0 17752 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698175906
transform 1 0 8736 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_171
timestamp 1698175906
transform 1 0 10248 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_201 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11928 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_158
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_162
timestamp 1698175906
transform 1 0 9744 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_192
timestamp 1698175906
transform 1 0 11424 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_196
timestamp 1698175906
transform 1 0 11648 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_204
timestamp 1698175906
transform 1 0 12096 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_152
timestamp 1698175906
transform 1 0 9184 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_156
timestamp 1698175906
transform 1 0 9408 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 10304 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 10416 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_183
timestamp 1698175906
transform 1 0 10920 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_187
timestamp 1698175906
transform 1 0 11144 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_218
timestamp 1698175906
transform 1 0 12880 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_222
timestamp 1698175906
transform 1 0 13104 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_238
timestamp 1698175906
transform 1 0 14000 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 14224 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698175906
transform 1 0 6720 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_110
timestamp 1698175906
transform 1 0 6832 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_153
timestamp 1698175906
transform 1 0 9240 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_191
timestamp 1698175906
transform 1 0 11368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_195
timestamp 1698175906
transform 1 0 11592 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_204
timestamp 1698175906
transform 1 0 12096 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_241
timestamp 1698175906
transform 1 0 14168 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_245
timestamp 1698175906
transform 1 0 14392 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_123
timestamp 1698175906
transform 1 0 7560 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_131
timestamp 1698175906
transform 1 0 8008 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_143
timestamp 1698175906
transform 1 0 8680 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_182
timestamp 1698175906
transform 1 0 10864 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_186
timestamp 1698175906
transform 1 0 11088 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_202
timestamp 1698175906
transform 1 0 11984 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_220
timestamp 1698175906
transform 1 0 12992 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_236
timestamp 1698175906
transform 1 0 13888 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 5152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_113
timestamp 1698175906
transform 1 0 7000 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_117
timestamp 1698175906
transform 1 0 7224 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_119
timestamp 1698175906
transform 1 0 7336 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_126
timestamp 1698175906
transform 1 0 7728 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_130
timestamp 1698175906
transform 1 0 7952 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_152
timestamp 1698175906
transform 1 0 9184 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_156
timestamp 1698175906
transform 1 0 9408 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_164
timestamp 1698175906
transform 1 0 9856 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_166
timestamp 1698175906
transform 1 0 9968 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_176
timestamp 1698175906
transform 1 0 10528 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_192
timestamp 1698175906
transform 1 0 11424 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_202
timestamp 1698175906
transform 1 0 11984 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 16128 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 4536 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698175906
transform 1 0 5432 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_93
timestamp 1698175906
transform 1 0 5880 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_120
timestamp 1698175906
transform 1 0 7392 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_152
timestamp 1698175906
transform 1 0 9184 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_160
timestamp 1698175906
transform 1 0 9632 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_169
timestamp 1698175906
transform 1 0 10136 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 10360 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_182
timestamp 1698175906
transform 1 0 10864 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_188
timestamp 1698175906
transform 1 0 11200 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_204
timestamp 1698175906
transform 1 0 12096 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_212
timestamp 1698175906
transform 1 0 12544 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_253
timestamp 1698175906
transform 1 0 14840 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_285
timestamp 1698175906
transform 1 0 16632 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_301
timestamp 1698175906
transform 1 0 17528 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_309
timestamp 1698175906
transform 1 0 17976 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698175906
transform 1 0 18200 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_92
timestamp 1698175906
transform 1 0 5824 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_118
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_134
timestamp 1698175906
transform 1 0 8176 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_177
timestamp 1698175906
transform 1 0 10584 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_179
timestamp 1698175906
transform 1 0 10696 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_185
timestamp 1698175906
transform 1 0 11032 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_195
timestamp 1698175906
transform 1 0 11592 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 12040 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_207
timestamp 1698175906
transform 1 0 12264 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_228
timestamp 1698175906
transform 1 0 13440 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_260
timestamp 1698175906
transform 1 0 15232 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 16128 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 4760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698175906
transform 1 0 6496 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_119
timestamp 1698175906
transform 1 0 7336 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698175906
transform 1 0 7784 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_129
timestamp 1698175906
transform 1 0 7896 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_141
timestamp 1698175906
transform 1 0 8568 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_151
timestamp 1698175906
transform 1 0 9128 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_158
timestamp 1698175906
transform 1 0 9520 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_195
timestamp 1698175906
transform 1 0 11592 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_212
timestamp 1698175906
transform 1 0 12544 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_106
timestamp 1698175906
transform 1 0 6608 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_135
timestamp 1698175906
transform 1 0 8232 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 8456 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_158
timestamp 1698175906
transform 1 0 9520 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_160
timestamp 1698175906
transform 1 0 9632 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_200
timestamp 1698175906
transform 1 0 11872 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698175906
transform 1 0 12656 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_244
timestamp 1698175906
transform 1 0 14336 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 16128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_111
timestamp 1698175906
transform 1 0 6888 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698175906
transform 1 0 10304 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 10416 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698175906
transform 1 0 10696 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_230
timestamp 1698175906
transform 1 0 13552 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_238
timestamp 1698175906
transform 1 0 14000 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 14224 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_96
timestamp 1698175906
transform 1 0 6048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_98
timestamp 1698175906
transform 1 0 6160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_128
timestamp 1698175906
transform 1 0 7840 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_198
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_225
timestamp 1698175906
transform 1 0 13272 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_257
timestamp 1698175906
transform 1 0 15064 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698175906
transform 1 0 15960 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 16184 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_120
timestamp 1698175906
transform 1 0 7392 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_138
timestamp 1698175906
transform 1 0 8400 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_142
timestamp 1698175906
transform 1 0 8624 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_190
timestamp 1698175906
transform 1 0 11312 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1698175906
transform 1 0 6496 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_117
timestamp 1698175906
transform 1 0 7224 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698175906
transform 1 0 8120 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_156
timestamp 1698175906
transform 1 0 9408 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_160
timestamp 1698175906
transform 1 0 9632 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_162
timestamp 1698175906
transform 1 0 9744 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_168
timestamp 1698175906
transform 1 0 10080 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_170
timestamp 1698175906
transform 1 0 10192 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_177
timestamp 1698175906
transform 1 0 10584 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_185
timestamp 1698175906
transform 1 0 11032 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_189
timestamp 1698175906
transform 1 0 11256 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_216
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_118
timestamp 1698175906
transform 1 0 7280 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_159
timestamp 1698175906
transform 1 0 9576 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698175906
transform 1 0 9800 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 10248 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_184
timestamp 1698175906
transform 1 0 10976 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_192
timestamp 1698175906
transform 1 0 11424 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_229
timestamp 1698175906
transform 1 0 13496 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_233
timestamp 1698175906
transform 1 0 13720 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 5152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_84
timestamp 1698175906
transform 1 0 5376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_114
timestamp 1698175906
transform 1 0 7056 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_118
timestamp 1698175906
transform 1 0 7280 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698175906
transform 1 0 8176 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_153
timestamp 1698175906
transform 1 0 9240 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_161
timestamp 1698175906
transform 1 0 9688 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_191
timestamp 1698175906
transform 1 0 11368 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_195
timestamp 1698175906
transform 1 0 11592 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_199
timestamp 1698175906
transform 1 0 11816 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_247
timestamp 1698175906
transform 1 0 14504 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_251
timestamp 1698175906
transform 1 0 14728 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_267
timestamp 1698175906
transform 1 0 15624 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1698175906
transform 1 0 16072 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_69
timestamp 1698175906
transform 1 0 4536 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_73
timestamp 1698175906
transform 1 0 4760 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_75
timestamp 1698175906
transform 1 0 4872 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_111
timestamp 1698175906
transform 1 0 6888 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_115
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_127
timestamp 1698175906
transform 1 0 7784 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_135
timestamp 1698175906
transform 1 0 8232 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_147
timestamp 1698175906
transform 1 0 8904 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_163
timestamp 1698175906
transform 1 0 9800 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 10248 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_182
timestamp 1698175906
transform 1 0 10864 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_198
timestamp 1698175906
transform 1 0 11760 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_206
timestamp 1698175906
transform 1 0 12208 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_210
timestamp 1698175906
transform 1 0 12432 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_212
timestamp 1698175906
transform 1 0 12544 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_223
timestamp 1698175906
transform 1 0 13160 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_239
timestamp 1698175906
transform 1 0 14056 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 14280 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 6720 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 6832 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_146
timestamp 1698175906
transform 1 0 8848 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_150
timestamp 1698175906
transform 1 0 9072 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_156
timestamp 1698175906
transform 1 0 9408 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_164
timestamp 1698175906
transform 1 0 9856 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_174
timestamp 1698175906
transform 1 0 10416 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_190
timestamp 1698175906
transform 1 0 11312 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_204
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_131
timestamp 1698175906
transform 1 0 8008 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_135
timestamp 1698175906
transform 1 0 8232 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_168
timestamp 1698175906
transform 1 0 10080 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 10416 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_179
timestamp 1698175906
transform 1 0 10696 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_182
timestamp 1698175906
transform 1 0 10864 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_190
timestamp 1698175906
transform 1 0 11312 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_220
timestamp 1698175906
transform 1 0 12992 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_224
timestamp 1698175906
transform 1 0 13216 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_240
timestamp 1698175906
transform 1 0 14112 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_150
timestamp 1698175906
transform 1 0 9072 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_180
timestamp 1698175906
transform 1 0 10752 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_217
timestamp 1698175906
transform 1 0 12824 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_221
timestamp 1698175906
transform 1 0 13048 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_253
timestamp 1698175906
transform 1 0 14840 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_269
timestamp 1698175906
transform 1 0 15736 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_277
timestamp 1698175906
transform 1 0 16184 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 16296 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_139
timestamp 1698175906
transform 1 0 8456 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_155
timestamp 1698175906
transform 1 0 9352 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698175906
transform 1 0 10360 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_193
timestamp 1698175906
transform 1 0 11480 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_199
timestamp 1698175906
transform 1 0 11816 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_203
timestamp 1698175906
transform 1 0 12040 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_210
timestamp 1698175906
transform 1 0 12432 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 14336 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_209
timestamp 1698175906
transform 1 0 12376 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698175906
transform 1 0 14280 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_144
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_171
timestamp 1698175906
transform 1 0 10248 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 11928 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita24_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13888 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita24_26
timestamp 1698175906
transform -1 0 17416 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 10472 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 8792 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 8792 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 12488 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 10472 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 12824 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 13104 20600 13160 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 17136 0 17192 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 10752 400 10808 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 13244 9772 13244 9772 0 _000_
rlabel metal2 6076 9072 6076 9072 0 _001_
rlabel metal2 7252 10570 7252 10570 0 _002_
rlabel metal3 7000 9940 7000 9940 0 _003_
rlabel metal2 12908 10248 12908 10248 0 _004_
rlabel metal2 9604 14196 9604 14196 0 _005_
rlabel metal2 11732 7420 11732 7420 0 _006_
rlabel metal2 6412 12376 6412 12376 0 _007_
rlabel metal2 9156 13342 9156 13342 0 _008_
rlabel metal2 6580 12516 6580 12516 0 _009_
rlabel metal2 10976 6916 10976 6916 0 _010_
rlabel metal2 7364 8008 7364 8008 0 _011_
rlabel metal3 8960 11900 8960 11900 0 _012_
rlabel metal2 11284 14196 11284 14196 0 _013_
rlabel metal3 12712 12292 12712 12292 0 _014_
rlabel metal2 12320 11508 12320 11508 0 _015_
rlabel metal2 7364 12880 7364 12880 0 _016_
rlabel metal2 13272 8876 13272 8876 0 _017_
rlabel metal2 12572 11200 12572 11200 0 _018_
rlabel metal2 8036 7434 8036 7434 0 _019_
rlabel metal2 13020 7812 13020 7812 0 _020_
rlabel metal2 10892 12152 10892 12152 0 _021_
rlabel metal3 10024 7700 10024 7700 0 _022_
rlabel metal2 6076 10696 6076 10696 0 _023_
rlabel metal2 11844 13356 11844 13356 0 _024_
rlabel metal2 7196 11200 7196 11200 0 _025_
rlabel metal2 6916 11984 6916 11984 0 _026_
rlabel metal2 9324 12068 9324 12068 0 _027_
rlabel metal3 9716 14196 9716 14196 0 _028_
rlabel metal2 6916 11676 6916 11676 0 _029_
rlabel metal2 10724 7224 10724 7224 0 _030_
rlabel metal2 10892 7406 10892 7406 0 _031_
rlabel metal2 8316 8820 8316 8820 0 _032_
rlabel metal2 9492 11340 9492 11340 0 _033_
rlabel metal2 8204 8400 8204 8400 0 _034_
rlabel metal2 9156 9548 9156 9548 0 _035_
rlabel metal2 8120 8484 8120 8484 0 _036_
rlabel metal2 9156 11816 9156 11816 0 _037_
rlabel metal3 9940 11900 9940 11900 0 _038_
rlabel metal2 11788 11816 11788 11816 0 _039_
rlabel metal2 11564 13342 11564 13342 0 _040_
rlabel metal2 12236 11956 12236 11956 0 _041_
rlabel metal2 12236 12544 12236 12544 0 _042_
rlabel metal2 11564 11788 11564 11788 0 _043_
rlabel metal2 10808 11844 10808 11844 0 _044_
rlabel metal2 12012 11704 12012 11704 0 _045_
rlabel metal3 10976 11564 10976 11564 0 _046_
rlabel metal2 12124 11844 12124 11844 0 _047_
rlabel metal2 9044 12488 9044 12488 0 _048_
rlabel metal2 8820 9912 8820 9912 0 _049_
rlabel metal3 8428 12460 8428 12460 0 _050_
rlabel metal2 11620 8512 11620 8512 0 _051_
rlabel metal2 10892 9128 10892 9128 0 _052_
rlabel metal2 10612 8624 10612 8624 0 _053_
rlabel metal2 11060 9100 11060 9100 0 _054_
rlabel metal2 13188 9212 13188 9212 0 _055_
rlabel metal2 13244 10920 13244 10920 0 _056_
rlabel metal2 8652 7896 8652 7896 0 _057_
rlabel metal3 12600 8036 12600 8036 0 _058_
rlabel metal2 10724 11956 10724 11956 0 _059_
rlabel metal3 11004 8428 11004 8428 0 _060_
rlabel metal2 10612 8232 10612 8232 0 _061_
rlabel metal3 7028 11116 7028 11116 0 _062_
rlabel metal3 9800 9996 9800 9996 0 _063_
rlabel metal3 9324 9940 9324 9940 0 _064_
rlabel metal3 8400 10052 8400 10052 0 _065_
rlabel metal2 8484 9660 8484 9660 0 _066_
rlabel metal2 6748 11284 6748 11284 0 _067_
rlabel metal2 6748 9352 6748 9352 0 _068_
rlabel metal2 6468 9184 6468 9184 0 _069_
rlabel metal3 7252 10052 7252 10052 0 _070_
rlabel metal2 8792 10780 8792 10780 0 _071_
rlabel metal2 11284 11116 11284 11116 0 _072_
rlabel metal2 10276 10584 10276 10584 0 _073_
rlabel metal2 6916 9940 6916 9940 0 _074_
rlabel metal2 6972 10612 6972 10612 0 _075_
rlabel metal2 7420 11340 7420 11340 0 _076_
rlabel metal2 12012 10612 12012 10612 0 _077_
rlabel metal3 11816 11956 11816 11956 0 _078_
rlabel metal2 6916 11816 6916 11816 0 _079_
rlabel metal3 11032 13244 11032 13244 0 _080_
rlabel metal3 12348 13804 12348 13804 0 _081_
rlabel metal2 11116 10556 11116 10556 0 _082_
rlabel metal2 11060 11228 11060 11228 0 _083_
rlabel metal2 12376 9996 12376 9996 0 _084_
rlabel metal2 12348 7728 12348 7728 0 _085_
rlabel metal2 8932 10220 8932 10220 0 _086_
rlabel metal2 11256 9660 11256 9660 0 _087_
rlabel metal2 10388 9324 10388 9324 0 _088_
rlabel metal2 9884 9604 9884 9604 0 _089_
rlabel metal2 10500 9240 10500 9240 0 _090_
rlabel metal2 12068 9772 12068 9772 0 _091_
rlabel metal2 7280 9548 7280 9548 0 _092_
rlabel metal2 8036 9772 8036 9772 0 _093_
rlabel metal2 12348 9464 12348 9464 0 _094_
rlabel metal2 12460 10164 12460 10164 0 _095_
rlabel metal2 9772 8624 9772 8624 0 _096_
rlabel metal2 9884 11536 9884 11536 0 _097_
rlabel metal2 10164 13916 10164 13916 0 _098_
rlabel metal2 11900 7728 11900 7728 0 _099_
rlabel metal3 9688 11508 9688 11508 0 _100_
rlabel metal2 11172 8540 11172 8540 0 _101_
rlabel metal2 11788 8400 11788 8400 0 _102_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal2 10836 10556 10836 10556 0 clknet_0_clk
rlabel metal2 6468 10416 6468 10416 0 clknet_1_0__leaf_clk
rlabel metal2 14644 12124 14644 12124 0 clknet_1_1__leaf_clk
rlabel metal2 6916 8428 6916 8428 0 dut24.count\[0\]
rlabel metal2 7028 9044 7028 9044 0 dut24.count\[1\]
rlabel metal2 8120 11172 8120 11172 0 dut24.count\[2\]
rlabel metal2 11284 9968 11284 9968 0 dut24.count\[3\]
rlabel metal2 13020 12908 13020 12908 0 net1
rlabel metal2 14084 12320 14084 12320 0 net10
rlabel metal2 10724 12460 10724 12460 0 net11
rlabel metal2 8484 4228 8484 4228 0 net12
rlabel metal2 10724 2982 10724 2982 0 net13
rlabel metal2 9100 6860 9100 6860 0 net14
rlabel metal2 14084 7616 14084 7616 0 net15
rlabel metal3 3178 12348 3178 12348 0 net16
rlabel metal3 10024 14252 10024 14252 0 net17
rlabel metal3 3178 12740 3178 12740 0 net18
rlabel metal2 12628 2982 12628 2982 0 net19
rlabel metal2 10556 3178 10556 3178 0 net2
rlabel metal2 10668 16240 10668 16240 0 net20
rlabel metal2 14308 9632 14308 9632 0 net21
rlabel metal2 12684 16128 12684 16128 0 net22
rlabel metal2 12348 14672 12348 14672 0 net23
rlabel metal2 5012 10808 5012 10808 0 net24
rlabel metal2 13132 19789 13132 19789 0 net25
rlabel metal2 17164 1015 17164 1015 0 net26
rlabel metal2 14252 11060 14252 11060 0 net3
rlabel metal2 8540 12936 8540 12936 0 net4
rlabel metal2 18956 8960 18956 8960 0 net5
rlabel metal3 3178 11956 3178 11956 0 net6
rlabel metal2 14644 8848 14644 8848 0 net7
rlabel metal2 12236 16660 12236 16660 0 net8
rlabel metal3 15190 12404 15190 12404 0 net9
rlabel metal2 19964 12936 19964 12936 0 segm[10]
rlabel metal2 10444 1211 10444 1211 0 segm[11]
rlabel metal2 20020 11004 20020 11004 0 segm[12]
rlabel metal3 9072 18732 9072 18732 0 segm[13]
rlabel metal3 20321 9100 20321 9100 0 segm[1]
rlabel metal3 679 11788 679 11788 0 segm[2]
rlabel metal2 20020 8820 20020 8820 0 segm[4]
rlabel metal3 12460 19124 12460 19124 0 segm[5]
rlabel metal2 20020 12628 20020 12628 0 segm[6]
rlabel metal2 20020 12180 20020 12180 0 segm[7]
rlabel metal2 11116 19971 11116 19971 0 segm[8]
rlabel metal2 8764 1211 8764 1211 0 segm[9]
rlabel metal2 11116 1015 11116 1015 0 sel[0]
rlabel metal2 9100 1099 9100 1099 0 sel[10]
rlabel metal2 20020 7924 20020 7924 0 sel[11]
rlabel metal3 679 12124 679 12124 0 sel[1]
rlabel metal2 9772 19971 9772 19971 0 sel[2]
rlabel metal3 679 12460 679 12460 0 sel[3]
rlabel metal2 12460 1099 12460 1099 0 sel[4]
rlabel metal3 10752 18732 10752 18732 0 sel[5]
rlabel metal2 20020 9548 20020 9548 0 sel[6]
rlabel metal2 12796 20573 12796 20573 0 sel[7]
rlabel metal3 12796 18732 12796 18732 0 sel[8]
rlabel metal3 679 10780 679 10780 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
