magic
tech gf180mcuD
magscale 1 5
timestamp 1699642761
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9417 19055 9423 19081
rect 9449 19055 9455 19081
rect 9865 18999 9871 19025
rect 9897 18999 9903 19025
rect 10705 18999 10711 19025
rect 10737 18999 10743 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 11047 18745 11073 18751
rect 11047 18713 11073 18719
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 10537 18607 10543 18633
rect 10569 18607 10575 18633
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 9535 13257 9561 13263
rect 9535 13225 9561 13231
rect 10263 13257 10289 13263
rect 10263 13225 10289 13231
rect 11383 13257 11409 13263
rect 11383 13225 11409 13231
rect 9591 13145 9617 13151
rect 9591 13113 9617 13119
rect 10319 13145 10345 13151
rect 10319 13113 10345 13119
rect 10823 13145 10849 13151
rect 10823 13113 10849 13119
rect 10935 13145 10961 13151
rect 10935 13113 10961 13119
rect 11159 13145 11185 13151
rect 11159 13113 11185 13119
rect 11271 13145 11297 13151
rect 11271 13113 11297 13119
rect 11439 13145 11465 13151
rect 11439 13113 11465 13119
rect 10879 13089 10905 13095
rect 10879 13057 10905 13063
rect 9535 13033 9561 13039
rect 9535 13001 9561 13007
rect 10263 13033 10289 13039
rect 10263 13001 10289 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 10313 12783 10319 12809
rect 10345 12783 10351 12809
rect 12329 12783 12335 12809
rect 12361 12783 12367 12809
rect 8857 12727 8863 12753
rect 8889 12727 8895 12753
rect 10929 12727 10935 12753
rect 10961 12727 10967 12753
rect 8247 12697 8273 12703
rect 13231 12697 13257 12703
rect 9249 12671 9255 12697
rect 9281 12671 9287 12697
rect 11265 12671 11271 12697
rect 11297 12671 11303 12697
rect 8247 12665 8273 12671
rect 13231 12665 13257 12671
rect 8079 12641 8105 12647
rect 8079 12609 8105 12615
rect 8191 12641 8217 12647
rect 8191 12609 8217 12615
rect 13063 12641 13089 12647
rect 13063 12609 13089 12615
rect 13175 12641 13201 12647
rect 13175 12609 13201 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 9535 12473 9561 12479
rect 9535 12441 9561 12447
rect 11999 12473 12025 12479
rect 11999 12441 12025 12447
rect 12055 12417 12081 12423
rect 7233 12391 7239 12417
rect 7265 12391 7271 12417
rect 10705 12391 10711 12417
rect 10737 12391 10743 12417
rect 12055 12385 12081 12391
rect 8807 12361 8833 12367
rect 6897 12335 6903 12361
rect 6929 12335 6935 12361
rect 8807 12329 8833 12335
rect 8919 12361 8945 12367
rect 9479 12361 9505 12367
rect 9081 12335 9087 12361
rect 9113 12335 9119 12361
rect 8919 12329 8945 12335
rect 9479 12329 9505 12335
rect 9591 12361 9617 12367
rect 9591 12329 9617 12335
rect 9815 12361 9841 12367
rect 11887 12361 11913 12367
rect 10369 12335 10375 12361
rect 10401 12335 10407 12361
rect 12609 12335 12615 12361
rect 12641 12335 12647 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 9815 12329 9841 12335
rect 11887 12329 11913 12335
rect 8863 12305 8889 12311
rect 8297 12279 8303 12305
rect 8329 12279 8335 12305
rect 11769 12279 11775 12305
rect 11801 12279 11807 12305
rect 13001 12279 13007 12305
rect 13033 12279 13039 12305
rect 14065 12279 14071 12305
rect 14097 12279 14103 12305
rect 8863 12273 8889 12279
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 11327 12025 11353 12031
rect 8465 11999 8471 12025
rect 8497 11999 8503 12025
rect 9529 11999 9535 12025
rect 9561 11999 9567 12025
rect 11327 11993 11353 11999
rect 12223 12025 12249 12031
rect 20007 12025 20033 12031
rect 14065 11999 14071 12025
rect 14097 11999 14103 12025
rect 12223 11993 12249 11999
rect 20007 11993 20033 11999
rect 11607 11969 11633 11975
rect 8129 11943 8135 11969
rect 8161 11943 8167 11969
rect 11607 11937 11633 11943
rect 12503 11969 12529 11975
rect 12609 11943 12615 11969
rect 12641 11943 12647 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 12503 11937 12529 11943
rect 11271 11913 11297 11919
rect 13001 11887 13007 11913
rect 13033 11887 13039 11913
rect 11271 11881 11297 11887
rect 11383 11857 11409 11863
rect 11383 11825 11409 11831
rect 12167 11857 12193 11863
rect 12167 11825 12193 11831
rect 12279 11857 12305 11863
rect 12279 11825 12305 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 8415 11689 8441 11695
rect 12671 11689 12697 11695
rect 9921 11663 9927 11689
rect 9953 11663 9959 11689
rect 10537 11663 10543 11689
rect 10569 11663 10575 11689
rect 8415 11657 8441 11663
rect 12671 11657 12697 11663
rect 12727 11689 12753 11695
rect 12727 11657 12753 11663
rect 13287 11689 13313 11695
rect 13287 11657 13313 11663
rect 8303 11633 8329 11639
rect 8303 11601 8329 11607
rect 8695 11633 8721 11639
rect 8695 11601 8721 11607
rect 13231 11633 13257 11639
rect 13231 11601 13257 11607
rect 8247 11577 8273 11583
rect 10711 11577 10737 11583
rect 10033 11551 10039 11577
rect 10065 11551 10071 11577
rect 8247 11545 8273 11551
rect 10711 11545 10737 11551
rect 12783 11577 12809 11583
rect 12783 11545 12809 11551
rect 13007 11577 13033 11583
rect 13007 11545 13033 11551
rect 8751 11465 8777 11471
rect 8751 11433 8777 11439
rect 13287 11465 13313 11471
rect 13287 11433 13313 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 7401 11215 7407 11241
rect 7433 11215 7439 11241
rect 8129 11215 8135 11241
rect 8161 11215 8167 11241
rect 7687 11185 7713 11191
rect 8639 11185 8665 11191
rect 7457 11159 7463 11185
rect 7489 11159 7495 11185
rect 8185 11159 8191 11185
rect 8217 11159 8223 11185
rect 7687 11153 7713 11159
rect 8639 11153 8665 11159
rect 8919 11185 8945 11191
rect 8919 11153 8945 11159
rect 9871 11185 9897 11191
rect 9871 11153 9897 11159
rect 10151 11185 10177 11191
rect 10151 11153 10177 11159
rect 10599 11185 10625 11191
rect 10599 11153 10625 11159
rect 8975 11129 9001 11135
rect 8129 11103 8135 11129
rect 8161 11103 8167 11129
rect 8975 11097 9001 11103
rect 10711 11129 10737 11135
rect 10711 11097 10737 11103
rect 10767 11129 10793 11135
rect 11153 11103 11159 11129
rect 11185 11103 11191 11129
rect 10767 11097 10793 11103
rect 7855 11073 7881 11079
rect 7855 11041 7881 11047
rect 8695 11073 8721 11079
rect 8695 11041 8721 11047
rect 8807 11073 8833 11079
rect 8807 11041 8833 11047
rect 9087 11073 9113 11079
rect 9087 11041 9113 11047
rect 9815 11073 9841 11079
rect 9815 11041 9841 11047
rect 9927 11073 9953 11079
rect 9927 11041 9953 11047
rect 10991 11073 11017 11079
rect 10991 11041 11017 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8023 10905 8049 10911
rect 8023 10873 8049 10879
rect 8135 10905 8161 10911
rect 8135 10873 8161 10879
rect 13063 10849 13089 10855
rect 7233 10823 7239 10849
rect 7265 10823 7271 10849
rect 9641 10823 9647 10849
rect 9673 10823 9679 10849
rect 13063 10817 13089 10823
rect 13455 10849 13481 10855
rect 13455 10817 13481 10823
rect 13511 10849 13537 10855
rect 13511 10817 13537 10823
rect 8303 10793 8329 10799
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 7625 10767 7631 10793
rect 7657 10767 7663 10793
rect 8303 10761 8329 10767
rect 8695 10793 8721 10799
rect 8695 10761 8721 10767
rect 8807 10793 8833 10799
rect 13119 10793 13145 10799
rect 9305 10767 9311 10793
rect 9337 10767 9343 10793
rect 10929 10767 10935 10793
rect 10961 10767 10967 10793
rect 8807 10761 8833 10767
rect 13119 10761 13145 10767
rect 13343 10793 13369 10799
rect 18937 10767 18943 10793
rect 18969 10767 18975 10793
rect 13343 10761 13369 10767
rect 6169 10711 6175 10737
rect 6201 10711 6207 10737
rect 10705 10711 10711 10737
rect 10737 10711 10743 10737
rect 11265 10711 11271 10737
rect 11297 10711 11303 10737
rect 12329 10711 12335 10737
rect 12361 10711 12367 10737
rect 19945 10711 19951 10737
rect 19977 10711 19983 10737
rect 967 10681 993 10687
rect 967 10649 993 10655
rect 7967 10681 7993 10687
rect 13063 10681 13089 10687
rect 8969 10655 8975 10681
rect 9001 10655 9007 10681
rect 7967 10649 7993 10655
rect 13063 10649 13089 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 14183 10513 14209 10519
rect 14183 10481 14209 10487
rect 7463 10457 7489 10463
rect 7463 10425 7489 10431
rect 10823 10457 10849 10463
rect 10823 10425 10849 10431
rect 20007 10457 20033 10463
rect 20007 10425 20033 10431
rect 6903 10401 6929 10407
rect 6903 10369 6929 10375
rect 6959 10401 6985 10407
rect 6959 10369 6985 10375
rect 7071 10401 7097 10407
rect 7071 10369 7097 10375
rect 7351 10401 7377 10407
rect 10935 10401 10961 10407
rect 14127 10401 14153 10407
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 11321 10375 11327 10401
rect 11353 10375 11359 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 7351 10369 7377 10375
rect 10935 10369 10961 10375
rect 14127 10369 14153 10375
rect 7575 10345 7601 10351
rect 7233 10319 7239 10345
rect 7265 10319 7271 10345
rect 9361 10319 9367 10345
rect 9393 10319 9399 10345
rect 12721 10319 12727 10345
rect 12753 10319 12759 10345
rect 7575 10313 7601 10319
rect 7351 10289 7377 10295
rect 14183 10289 14209 10295
rect 11097 10263 11103 10289
rect 11129 10263 11135 10289
rect 7351 10257 7377 10263
rect 14183 10257 14209 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 7905 10095 7911 10121
rect 7937 10095 7943 10121
rect 7121 10039 7127 10065
rect 7153 10039 7159 10065
rect 8073 10039 8079 10065
rect 8105 10039 8111 10065
rect 8241 10039 8247 10065
rect 8273 10039 8279 10065
rect 11321 10039 11327 10065
rect 11353 10039 11359 10065
rect 13113 10039 13119 10065
rect 13145 10039 13151 10065
rect 9031 10009 9057 10015
rect 7513 9983 7519 10009
rect 7545 9983 7551 10009
rect 8353 9983 8359 10009
rect 8385 9983 8391 10009
rect 9417 9983 9423 10009
rect 9449 9983 9455 10009
rect 9641 9983 9647 10009
rect 9673 9983 9679 10009
rect 12721 9983 12727 10009
rect 12753 9983 12759 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 9031 9977 9057 9983
rect 6057 9927 6063 9953
rect 6089 9927 6095 9953
rect 9249 9927 9255 9953
rect 9281 9927 9287 9953
rect 14177 9927 14183 9953
rect 14209 9927 14215 9953
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 967 9673 993 9679
rect 967 9641 993 9647
rect 10767 9673 10793 9679
rect 10767 9641 10793 9647
rect 11663 9673 11689 9679
rect 11663 9641 11689 9647
rect 12111 9673 12137 9679
rect 12111 9641 12137 9647
rect 20007 9673 20033 9679
rect 20007 9641 20033 9647
rect 7799 9617 7825 9623
rect 2137 9591 2143 9617
rect 2169 9591 2175 9617
rect 7799 9585 7825 9591
rect 8191 9617 8217 9623
rect 8191 9585 8217 9591
rect 8359 9617 8385 9623
rect 8359 9585 8385 9591
rect 9311 9617 9337 9623
rect 9311 9585 9337 9591
rect 9983 9617 10009 9623
rect 9983 9585 10009 9591
rect 11551 9617 11577 9623
rect 11551 9585 11577 9591
rect 11775 9617 11801 9623
rect 12049 9591 12055 9617
rect 12081 9591 12087 9617
rect 12721 9591 12727 9617
rect 12753 9591 12759 9617
rect 14625 9591 14631 9617
rect 14657 9591 14663 9617
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 11775 9585 11801 9591
rect 7967 9561 7993 9567
rect 7967 9529 7993 9535
rect 8079 9561 8105 9567
rect 8079 9529 8105 9535
rect 8303 9561 8329 9567
rect 8303 9529 8329 9535
rect 9143 9561 9169 9567
rect 10823 9561 10849 9567
rect 9529 9535 9535 9561
rect 9561 9535 9567 9561
rect 9809 9535 9815 9561
rect 9841 9535 9847 9561
rect 9143 9529 9169 9535
rect 10823 9529 10849 9535
rect 10991 9561 11017 9567
rect 10991 9529 11017 9535
rect 11383 9561 11409 9567
rect 11383 9529 11409 9535
rect 11887 9561 11913 9567
rect 11887 9529 11913 9535
rect 12279 9561 12305 9567
rect 13113 9535 13119 9561
rect 13145 9535 13151 9561
rect 12279 9529 12305 9535
rect 7855 9505 7881 9511
rect 7855 9473 7881 9479
rect 9255 9505 9281 9511
rect 10375 9505 10401 9511
rect 9977 9479 9983 9505
rect 10009 9479 10015 9505
rect 10201 9479 10207 9505
rect 10233 9479 10239 9505
rect 9255 9473 9281 9479
rect 10375 9473 10401 9479
rect 10711 9505 10737 9511
rect 10711 9473 10737 9479
rect 11047 9505 11073 9511
rect 11047 9473 11073 9479
rect 11159 9505 11185 9511
rect 11159 9473 11185 9479
rect 11215 9505 11241 9511
rect 11215 9473 11241 9479
rect 11327 9505 11353 9511
rect 11327 9473 11353 9479
rect 12167 9505 12193 9511
rect 14233 9479 14239 9505
rect 14265 9479 14271 9505
rect 14737 9479 14743 9505
rect 14769 9479 14775 9505
rect 12167 9473 12193 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 11047 9337 11073 9343
rect 13231 9337 13257 9343
rect 8745 9311 8751 9337
rect 8777 9311 8783 9337
rect 10761 9311 10767 9337
rect 10793 9311 10799 9337
rect 12609 9311 12615 9337
rect 12641 9311 12647 9337
rect 11047 9305 11073 9311
rect 13231 9305 13257 9311
rect 9367 9281 9393 9287
rect 9367 9249 9393 9255
rect 9535 9281 9561 9287
rect 9535 9249 9561 9255
rect 9647 9281 9673 9287
rect 13343 9281 13369 9287
rect 10313 9255 10319 9281
rect 10345 9255 10351 9281
rect 9647 9249 9673 9255
rect 13343 9249 13369 9255
rect 13399 9281 13425 9287
rect 14457 9255 14463 9281
rect 14489 9255 14495 9281
rect 13399 9249 13425 9255
rect 8919 9225 8945 9231
rect 7289 9199 7295 9225
rect 7321 9199 7327 9225
rect 7681 9199 7687 9225
rect 7713 9199 7719 9225
rect 8919 9193 8945 9199
rect 9703 9225 9729 9231
rect 9703 9193 9729 9199
rect 9871 9225 9897 9231
rect 9871 9193 9897 9199
rect 10151 9225 10177 9231
rect 10593 9199 10599 9225
rect 10625 9199 10631 9225
rect 10873 9199 10879 9225
rect 10905 9199 10911 9225
rect 12721 9199 12727 9225
rect 12753 9199 12759 9225
rect 14345 9199 14351 9225
rect 14377 9199 14383 9225
rect 18937 9199 18943 9225
rect 18969 9199 18975 9225
rect 10151 9193 10177 9199
rect 9311 9169 9337 9175
rect 6225 9143 6231 9169
rect 6257 9143 6263 9169
rect 9311 9137 9337 9143
rect 11103 9169 11129 9175
rect 11103 9137 11129 9143
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 12559 8889 12585 8895
rect 12559 8857 12585 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 8359 8833 8385 8839
rect 9087 8833 9113 8839
rect 9479 8833 9505 8839
rect 8129 8807 8135 8833
rect 8161 8807 8167 8833
rect 8801 8807 8807 8833
rect 8833 8807 8839 8833
rect 9193 8807 9199 8833
rect 9225 8807 9231 8833
rect 8359 8801 8385 8807
rect 9087 8801 9113 8807
rect 9479 8801 9505 8807
rect 9591 8833 9617 8839
rect 9591 8801 9617 8807
rect 9759 8833 9785 8839
rect 9759 8801 9785 8807
rect 9927 8833 9953 8839
rect 9927 8801 9953 8807
rect 10823 8833 10849 8839
rect 10823 8801 10849 8807
rect 12055 8833 12081 8839
rect 12447 8833 12473 8839
rect 12329 8807 12335 8833
rect 12361 8807 12367 8833
rect 12609 8807 12615 8833
rect 12641 8807 12647 8833
rect 18937 8807 18943 8833
rect 18969 8807 18975 8833
rect 12055 8801 12081 8807
rect 12447 8801 12473 8807
rect 10095 8777 10121 8783
rect 10095 8745 10121 8751
rect 10207 8777 10233 8783
rect 10649 8751 10655 8777
rect 10681 8751 10687 8777
rect 10207 8745 10233 8751
rect 9703 8721 9729 8727
rect 8913 8695 8919 8721
rect 8945 8695 8951 8721
rect 9703 8689 9729 8695
rect 10151 8721 10177 8727
rect 10151 8689 10177 8695
rect 12111 8721 12137 8727
rect 12111 8689 12137 8695
rect 12167 8721 12193 8727
rect 12167 8689 12193 8695
rect 12727 8721 12753 8727
rect 12727 8689 12753 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 9703 8553 9729 8559
rect 9703 8521 9729 8527
rect 9815 8553 9841 8559
rect 9815 8521 9841 8527
rect 10207 8553 10233 8559
rect 10207 8521 10233 8527
rect 10319 8553 10345 8559
rect 10319 8521 10345 8527
rect 13119 8553 13145 8559
rect 13119 8521 13145 8527
rect 8751 8497 8777 8503
rect 7345 8471 7351 8497
rect 7377 8471 7383 8497
rect 8751 8465 8777 8471
rect 8863 8497 8889 8503
rect 8863 8465 8889 8471
rect 8975 8497 9001 8503
rect 8975 8465 9001 8471
rect 11887 8497 11913 8503
rect 13281 8471 13287 8497
rect 13313 8471 13319 8497
rect 11887 8465 11913 8471
rect 8639 8441 8665 8447
rect 10151 8441 10177 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 7009 8415 7015 8441
rect 7041 8415 7047 8441
rect 9977 8415 9983 8441
rect 10009 8415 10015 8441
rect 8639 8409 8665 8415
rect 10151 8409 10177 8415
rect 11495 8441 11521 8447
rect 11495 8409 11521 8415
rect 11607 8441 11633 8447
rect 11607 8409 11633 8415
rect 11775 8441 11801 8447
rect 11775 8409 11801 8415
rect 11999 8441 12025 8447
rect 11999 8409 12025 8415
rect 12223 8441 12249 8447
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 12223 8409 12249 8415
rect 9759 8385 9785 8391
rect 8409 8359 8415 8385
rect 8441 8359 8447 8385
rect 9759 8353 9785 8359
rect 11663 8385 11689 8391
rect 11663 8353 11689 8359
rect 12111 8385 12137 8391
rect 12111 8353 12137 8359
rect 20007 8385 20033 8391
rect 20007 8353 20033 8359
rect 967 8329 993 8335
rect 967 8297 993 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 9927 8105 9953 8111
rect 20007 8105 20033 8111
rect 7121 8079 7127 8105
rect 7153 8079 7159 8105
rect 8185 8079 8191 8105
rect 8217 8079 8223 8105
rect 12105 8079 12111 8105
rect 12137 8079 12143 8105
rect 13169 8079 13175 8105
rect 13201 8079 13207 8105
rect 9927 8073 9953 8079
rect 20007 8073 20033 8079
rect 8303 8049 8329 8055
rect 6785 8023 6791 8049
rect 6817 8023 6823 8049
rect 8303 8017 8329 8023
rect 8471 8049 8497 8055
rect 8471 8017 8497 8023
rect 9815 8049 9841 8055
rect 9815 8017 9841 8023
rect 10151 8049 10177 8055
rect 10151 8017 10177 8023
rect 10599 8049 10625 8055
rect 10599 8017 10625 8023
rect 10767 8049 10793 8055
rect 10767 8017 10793 8023
rect 10935 8049 10961 8055
rect 11769 8023 11775 8049
rect 11801 8023 11807 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 10935 8017 10961 8023
rect 10095 7993 10121 7999
rect 10095 7961 10121 7967
rect 8415 7937 8441 7943
rect 8415 7905 8441 7911
rect 10039 7937 10065 7943
rect 10039 7905 10065 7911
rect 10711 7937 10737 7943
rect 10711 7905 10737 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 7295 7769 7321 7775
rect 7295 7737 7321 7743
rect 10991 7769 11017 7775
rect 10991 7737 11017 7743
rect 12783 7769 12809 7775
rect 12783 7737 12809 7743
rect 7457 7687 7463 7713
rect 7489 7687 7495 7713
rect 7625 7687 7631 7713
rect 7657 7687 7663 7713
rect 8129 7687 8135 7713
rect 8161 7687 8167 7713
rect 9585 7687 9591 7713
rect 9617 7687 9623 7713
rect 10817 7687 10823 7713
rect 10849 7687 10855 7713
rect 12945 7687 12951 7713
rect 12977 7687 12983 7713
rect 7799 7657 7825 7663
rect 8017 7631 8023 7657
rect 8049 7631 8055 7657
rect 9249 7631 9255 7657
rect 9281 7631 9287 7657
rect 7799 7625 7825 7631
rect 10649 7575 10655 7601
rect 10681 7575 10687 7601
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 12049 7295 12055 7321
rect 12081 7295 12087 7321
rect 13113 7295 13119 7321
rect 13145 7295 13151 7321
rect 11713 7239 11719 7265
rect 11745 7239 11751 7265
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 10593 6903 10599 6929
rect 10625 6903 10631 6929
rect 10929 6847 10935 6873
rect 10961 6847 10967 6873
rect 9529 6791 9535 6817
rect 9561 6791 9567 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 8359 2617 8385 2623
rect 8359 2585 8385 2591
rect 7849 2535 7855 2561
rect 7881 2535 7887 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 10201 2143 10207 2169
rect 10233 2143 10239 2169
rect 10711 2057 10737 2063
rect 10711 2025 10737 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 11215 1833 11241 1839
rect 11215 1801 11241 1807
rect 13063 1833 13089 1839
rect 13063 1801 13089 1807
rect 7961 1751 7967 1777
rect 7993 1751 7999 1777
rect 8465 1751 8471 1777
rect 8497 1751 8503 1777
rect 10817 1751 10823 1777
rect 10849 1751 10855 1777
rect 12609 1751 12615 1777
rect 12641 1751 12647 1777
rect 7401 1695 7407 1721
rect 7433 1695 7439 1721
rect 9249 1695 9255 1721
rect 9281 1695 9287 1721
rect 4159 1665 4185 1671
rect 4159 1633 4185 1639
rect 15247 1665 15273 1671
rect 15247 1633 15273 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 9423 19055 9449 19081
rect 9871 18999 9897 19025
rect 10711 18999 10737 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 11047 18719 11073 18745
rect 13119 18719 13145 18745
rect 10543 18607 10569 18633
rect 12615 18607 12641 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 9535 13231 9561 13257
rect 10263 13231 10289 13257
rect 11383 13231 11409 13257
rect 9591 13119 9617 13145
rect 10319 13119 10345 13145
rect 10823 13119 10849 13145
rect 10935 13119 10961 13145
rect 11159 13119 11185 13145
rect 11271 13119 11297 13145
rect 11439 13119 11465 13145
rect 10879 13063 10905 13089
rect 9535 13007 9561 13033
rect 10263 13007 10289 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 10319 12783 10345 12809
rect 12335 12783 12361 12809
rect 8863 12727 8889 12753
rect 10935 12727 10961 12753
rect 8247 12671 8273 12697
rect 9255 12671 9281 12697
rect 11271 12671 11297 12697
rect 13231 12671 13257 12697
rect 8079 12615 8105 12641
rect 8191 12615 8217 12641
rect 13063 12615 13089 12641
rect 13175 12615 13201 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 9535 12447 9561 12473
rect 11999 12447 12025 12473
rect 7239 12391 7265 12417
rect 10711 12391 10737 12417
rect 12055 12391 12081 12417
rect 6903 12335 6929 12361
rect 8807 12335 8833 12361
rect 8919 12335 8945 12361
rect 9087 12335 9113 12361
rect 9479 12335 9505 12361
rect 9591 12335 9617 12361
rect 9815 12335 9841 12361
rect 10375 12335 10401 12361
rect 11887 12335 11913 12361
rect 12615 12335 12641 12361
rect 18831 12335 18857 12361
rect 8303 12279 8329 12305
rect 8863 12279 8889 12305
rect 11775 12279 11801 12305
rect 13007 12279 13033 12305
rect 14071 12279 14097 12305
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 8471 11999 8497 12025
rect 9535 11999 9561 12025
rect 11327 11999 11353 12025
rect 12223 11999 12249 12025
rect 14071 11999 14097 12025
rect 20007 11999 20033 12025
rect 8135 11943 8161 11969
rect 11607 11943 11633 11969
rect 12503 11943 12529 11969
rect 12615 11943 12641 11969
rect 18831 11943 18857 11969
rect 11271 11887 11297 11913
rect 13007 11887 13033 11913
rect 11383 11831 11409 11857
rect 12167 11831 12193 11857
rect 12279 11831 12305 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 8415 11663 8441 11689
rect 9927 11663 9953 11689
rect 10543 11663 10569 11689
rect 12671 11663 12697 11689
rect 12727 11663 12753 11689
rect 13287 11663 13313 11689
rect 8303 11607 8329 11633
rect 8695 11607 8721 11633
rect 13231 11607 13257 11633
rect 8247 11551 8273 11577
rect 10039 11551 10065 11577
rect 10711 11551 10737 11577
rect 12783 11551 12809 11577
rect 13007 11551 13033 11577
rect 8751 11439 8777 11465
rect 13287 11439 13313 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7407 11215 7433 11241
rect 8135 11215 8161 11241
rect 7463 11159 7489 11185
rect 7687 11159 7713 11185
rect 8191 11159 8217 11185
rect 8639 11159 8665 11185
rect 8919 11159 8945 11185
rect 9871 11159 9897 11185
rect 10151 11159 10177 11185
rect 10599 11159 10625 11185
rect 8135 11103 8161 11129
rect 8975 11103 9001 11129
rect 10711 11103 10737 11129
rect 10767 11103 10793 11129
rect 11159 11103 11185 11129
rect 7855 11047 7881 11073
rect 8695 11047 8721 11073
rect 8807 11047 8833 11073
rect 9087 11047 9113 11073
rect 9815 11047 9841 11073
rect 9927 11047 9953 11073
rect 10991 11047 11017 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8023 10879 8049 10905
rect 8135 10879 8161 10905
rect 7239 10823 7265 10849
rect 9647 10823 9673 10849
rect 13063 10823 13089 10849
rect 13455 10823 13481 10849
rect 13511 10823 13537 10849
rect 2143 10767 2169 10793
rect 7631 10767 7657 10793
rect 8303 10767 8329 10793
rect 8695 10767 8721 10793
rect 8807 10767 8833 10793
rect 9311 10767 9337 10793
rect 10935 10767 10961 10793
rect 13119 10767 13145 10793
rect 13343 10767 13369 10793
rect 18943 10767 18969 10793
rect 6175 10711 6201 10737
rect 10711 10711 10737 10737
rect 11271 10711 11297 10737
rect 12335 10711 12361 10737
rect 19951 10711 19977 10737
rect 967 10655 993 10681
rect 7967 10655 7993 10681
rect 8975 10655 9001 10681
rect 13063 10655 13089 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 14183 10487 14209 10513
rect 7463 10431 7489 10457
rect 10823 10431 10849 10457
rect 20007 10431 20033 10457
rect 6903 10375 6929 10401
rect 6959 10375 6985 10401
rect 7071 10375 7097 10401
rect 7351 10375 7377 10401
rect 10039 10375 10065 10401
rect 10935 10375 10961 10401
rect 11327 10375 11353 10401
rect 14127 10375 14153 10401
rect 18831 10375 18857 10401
rect 7239 10319 7265 10345
rect 7575 10319 7601 10345
rect 9367 10319 9393 10345
rect 12727 10319 12753 10345
rect 7351 10263 7377 10289
rect 11103 10263 11129 10289
rect 14183 10263 14209 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7911 10095 7937 10121
rect 7127 10039 7153 10065
rect 8079 10039 8105 10065
rect 8247 10039 8273 10065
rect 11327 10039 11353 10065
rect 13119 10039 13145 10065
rect 7519 9983 7545 10009
rect 8359 9983 8385 10009
rect 9031 9983 9057 10009
rect 9423 9983 9449 10009
rect 9647 9983 9673 10009
rect 12727 9983 12753 10009
rect 18831 9983 18857 10009
rect 6063 9927 6089 9953
rect 9255 9927 9281 9953
rect 14183 9927 14209 9953
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 967 9647 993 9673
rect 10767 9647 10793 9673
rect 11663 9647 11689 9673
rect 12111 9647 12137 9673
rect 20007 9647 20033 9673
rect 2143 9591 2169 9617
rect 7799 9591 7825 9617
rect 8191 9591 8217 9617
rect 8359 9591 8385 9617
rect 9311 9591 9337 9617
rect 9983 9591 10009 9617
rect 11551 9591 11577 9617
rect 11775 9591 11801 9617
rect 12055 9591 12081 9617
rect 12727 9591 12753 9617
rect 14631 9591 14657 9617
rect 18831 9591 18857 9617
rect 7967 9535 7993 9561
rect 8079 9535 8105 9561
rect 8303 9535 8329 9561
rect 9143 9535 9169 9561
rect 9535 9535 9561 9561
rect 9815 9535 9841 9561
rect 10823 9535 10849 9561
rect 10991 9535 11017 9561
rect 11383 9535 11409 9561
rect 11887 9535 11913 9561
rect 12279 9535 12305 9561
rect 13119 9535 13145 9561
rect 7855 9479 7881 9505
rect 9255 9479 9281 9505
rect 9983 9479 10009 9505
rect 10207 9479 10233 9505
rect 10375 9479 10401 9505
rect 10711 9479 10737 9505
rect 11047 9479 11073 9505
rect 11159 9479 11185 9505
rect 11215 9479 11241 9505
rect 11327 9479 11353 9505
rect 12167 9479 12193 9505
rect 14239 9479 14265 9505
rect 14743 9479 14769 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 8751 9311 8777 9337
rect 10767 9311 10793 9337
rect 11047 9311 11073 9337
rect 12615 9311 12641 9337
rect 13231 9311 13257 9337
rect 9367 9255 9393 9281
rect 9535 9255 9561 9281
rect 9647 9255 9673 9281
rect 10319 9255 10345 9281
rect 13343 9255 13369 9281
rect 13399 9255 13425 9281
rect 14463 9255 14489 9281
rect 7295 9199 7321 9225
rect 7687 9199 7713 9225
rect 8919 9199 8945 9225
rect 9703 9199 9729 9225
rect 9871 9199 9897 9225
rect 10151 9199 10177 9225
rect 10599 9199 10625 9225
rect 10879 9199 10905 9225
rect 12727 9199 12753 9225
rect 14351 9199 14377 9225
rect 18943 9199 18969 9225
rect 6231 9143 6257 9169
rect 9311 9143 9337 9169
rect 11103 9143 11129 9169
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 12559 8863 12585 8889
rect 20007 8863 20033 8889
rect 8135 8807 8161 8833
rect 8359 8807 8385 8833
rect 8807 8807 8833 8833
rect 9087 8807 9113 8833
rect 9199 8807 9225 8833
rect 9479 8807 9505 8833
rect 9591 8807 9617 8833
rect 9759 8807 9785 8833
rect 9927 8807 9953 8833
rect 10823 8807 10849 8833
rect 12055 8807 12081 8833
rect 12335 8807 12361 8833
rect 12447 8807 12473 8833
rect 12615 8807 12641 8833
rect 18943 8807 18969 8833
rect 10095 8751 10121 8777
rect 10207 8751 10233 8777
rect 10655 8751 10681 8777
rect 8919 8695 8945 8721
rect 9703 8695 9729 8721
rect 10151 8695 10177 8721
rect 12111 8695 12137 8721
rect 12167 8695 12193 8721
rect 12727 8695 12753 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 9703 8527 9729 8553
rect 9815 8527 9841 8553
rect 10207 8527 10233 8553
rect 10319 8527 10345 8553
rect 13119 8527 13145 8553
rect 7351 8471 7377 8497
rect 8751 8471 8777 8497
rect 8863 8471 8889 8497
rect 8975 8471 9001 8497
rect 11887 8471 11913 8497
rect 13287 8471 13313 8497
rect 2143 8415 2169 8441
rect 7015 8415 7041 8441
rect 8639 8415 8665 8441
rect 9983 8415 10009 8441
rect 10151 8415 10177 8441
rect 11495 8415 11521 8441
rect 11607 8415 11633 8441
rect 11775 8415 11801 8441
rect 11999 8415 12025 8441
rect 12223 8415 12249 8441
rect 18831 8415 18857 8441
rect 8415 8359 8441 8385
rect 9759 8359 9785 8385
rect 11663 8359 11689 8385
rect 12111 8359 12137 8385
rect 20007 8359 20033 8385
rect 967 8303 993 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 7127 8079 7153 8105
rect 8191 8079 8217 8105
rect 9927 8079 9953 8105
rect 12111 8079 12137 8105
rect 13175 8079 13201 8105
rect 20007 8079 20033 8105
rect 6791 8023 6817 8049
rect 8303 8023 8329 8049
rect 8471 8023 8497 8049
rect 9815 8023 9841 8049
rect 10151 8023 10177 8049
rect 10599 8023 10625 8049
rect 10767 8023 10793 8049
rect 10935 8023 10961 8049
rect 11775 8023 11801 8049
rect 18831 8023 18857 8049
rect 10095 7967 10121 7993
rect 8415 7911 8441 7937
rect 10039 7911 10065 7937
rect 10711 7911 10737 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 7295 7743 7321 7769
rect 10991 7743 11017 7769
rect 12783 7743 12809 7769
rect 7463 7687 7489 7713
rect 7631 7687 7657 7713
rect 8135 7687 8161 7713
rect 9591 7687 9617 7713
rect 10823 7687 10849 7713
rect 12951 7687 12977 7713
rect 7799 7631 7825 7657
rect 8023 7631 8049 7657
rect 9255 7631 9281 7657
rect 10655 7575 10681 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 12055 7295 12081 7321
rect 13119 7295 13145 7321
rect 11719 7239 11745 7265
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 10599 6903 10625 6929
rect 10935 6847 10961 6873
rect 9535 6791 9561 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 8359 2591 8385 2617
rect 7855 2535 7881 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 10207 2143 10233 2169
rect 10711 2031 10737 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 11215 1807 11241 1833
rect 13063 1807 13089 1833
rect 7967 1751 7993 1777
rect 8471 1751 8497 1777
rect 10823 1751 10849 1777
rect 12615 1751 12641 1777
rect 7407 1695 7433 1721
rect 9255 1695 9281 1721
rect 4159 1639 4185 1665
rect 15247 1639 15273 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 9408 20600 9464 21000
rect 10416 20600 10472 21000
rect 10752 20600 10808 21000
rect 11760 20600 11816 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 9422 19081 9450 20600
rect 9422 19055 9423 19081
rect 9449 19055 9450 19081
rect 9422 19049 9450 19055
rect 9870 19026 9898 19031
rect 9534 19025 9898 19026
rect 9534 18999 9871 19025
rect 9897 18999 9898 19025
rect 9534 18998 9898 18999
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 9534 13258 9562 18998
rect 9870 18993 9898 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10430 18746 10458 20600
rect 10766 19138 10794 20600
rect 10766 19105 10794 19110
rect 11214 19138 11242 19143
rect 11214 19091 11242 19110
rect 11774 19138 11802 20600
rect 11774 19105 11802 19110
rect 10430 18713 10458 18718
rect 10710 19025 10738 19031
rect 10710 18999 10711 19025
rect 10737 18999 10738 19025
rect 10542 18633 10570 18639
rect 10542 18607 10543 18633
rect 10569 18607 10570 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 10542 15974 10570 18607
rect 10710 15974 10738 18999
rect 11046 18746 11074 18751
rect 11046 18699 11074 18718
rect 12110 18746 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 12110 18713 12138 18718
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 10262 15946 10570 15974
rect 10654 15946 10738 15974
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10262 13258 10290 15946
rect 9534 13257 9674 13258
rect 9534 13231 9535 13257
rect 9561 13231 9674 13257
rect 9534 13230 9674 13231
rect 9534 13225 9562 13230
rect 9590 13145 9618 13151
rect 9590 13119 9591 13145
rect 9617 13119 9618 13145
rect 9086 13034 9114 13039
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2086 12810 2114 12815
rect 966 10681 994 10687
rect 966 10655 967 10681
rect 993 10655 994 10681
rect 966 10458 994 10655
rect 966 10425 994 10430
rect 2086 9954 2114 12782
rect 8862 12753 8890 12759
rect 8862 12727 8863 12753
rect 8889 12727 8890 12753
rect 8246 12698 8274 12703
rect 8246 12697 8386 12698
rect 8246 12671 8247 12697
rect 8273 12671 8386 12697
rect 8246 12670 8386 12671
rect 8246 12665 8274 12670
rect 7238 12642 7266 12647
rect 6902 12418 6930 12423
rect 6902 12361 6930 12390
rect 7238 12417 7266 12614
rect 8078 12642 8106 12647
rect 8078 12595 8106 12614
rect 8190 12642 8218 12647
rect 7238 12391 7239 12417
rect 7265 12391 7266 12417
rect 7238 12385 7266 12391
rect 7630 12418 7658 12423
rect 6902 12335 6903 12361
rect 6929 12335 6930 12361
rect 6902 12329 6930 12335
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 7406 11241 7434 11247
rect 7406 11215 7407 11241
rect 7433 11215 7434 11241
rect 6174 11186 6202 11191
rect 2142 10794 2170 10799
rect 2142 10747 2170 10766
rect 6062 10794 6090 10799
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2086 9921 2114 9926
rect 6062 10402 6090 10766
rect 6174 10737 6202 11158
rect 7406 11130 7434 11215
rect 7462 11186 7490 11205
rect 7462 11153 7490 11158
rect 7238 11102 7406 11130
rect 7238 10849 7266 11102
rect 7406 11097 7434 11102
rect 7238 10823 7239 10849
rect 7265 10823 7266 10849
rect 7238 10817 7266 10823
rect 7462 10962 7490 10967
rect 6174 10711 6175 10737
rect 6201 10711 6202 10737
rect 6174 10705 6202 10711
rect 7462 10457 7490 10934
rect 7630 10794 7658 12390
rect 8134 12418 8162 12423
rect 8134 11969 8162 12390
rect 8134 11943 8135 11969
rect 8161 11943 8162 11969
rect 8134 11937 8162 11943
rect 8190 11802 8218 12614
rect 8358 12362 8386 12670
rect 8862 12418 8890 12727
rect 8862 12385 8890 12390
rect 8134 11774 8218 11802
rect 8302 12305 8330 12311
rect 8302 12279 8303 12305
rect 8329 12279 8330 12305
rect 8134 11241 8162 11774
rect 8302 11746 8330 12279
rect 8134 11215 8135 11241
rect 8161 11215 8162 11241
rect 8134 11209 8162 11215
rect 8190 11718 8302 11746
rect 7686 11186 7714 11191
rect 7686 11139 7714 11158
rect 8190 11185 8218 11718
rect 8302 11713 8330 11718
rect 8358 11690 8386 12334
rect 8806 12362 8834 12367
rect 8806 12315 8834 12334
rect 8918 12361 8946 12367
rect 8918 12335 8919 12361
rect 8945 12335 8946 12361
rect 8862 12305 8890 12311
rect 8862 12279 8863 12305
rect 8889 12279 8890 12305
rect 8862 12138 8890 12279
rect 8918 12250 8946 12335
rect 9086 12361 9114 13006
rect 9534 13034 9562 13039
rect 9534 12987 9562 13006
rect 9254 12698 9282 12703
rect 9254 12697 9562 12698
rect 9254 12671 9255 12697
rect 9281 12671 9562 12697
rect 9254 12670 9562 12671
rect 9254 12665 9282 12670
rect 9534 12473 9562 12670
rect 9534 12447 9535 12473
rect 9561 12447 9562 12473
rect 9534 12441 9562 12447
rect 9590 12474 9618 13119
rect 9590 12441 9618 12446
rect 9086 12335 9087 12361
rect 9113 12335 9114 12361
rect 9086 12329 9114 12335
rect 9478 12361 9506 12367
rect 9478 12335 9479 12361
rect 9505 12335 9506 12361
rect 8918 12217 8946 12222
rect 8470 12110 8890 12138
rect 8470 12025 8498 12110
rect 8470 11999 8471 12025
rect 8497 11999 8498 12025
rect 8470 11993 8498 11999
rect 8694 11746 8722 11751
rect 8414 11690 8442 11695
rect 8358 11689 8442 11690
rect 8358 11663 8415 11689
rect 8441 11663 8442 11689
rect 8358 11662 8442 11663
rect 8414 11657 8442 11662
rect 8302 11634 8330 11639
rect 8694 11634 8722 11718
rect 8302 11633 8386 11634
rect 8302 11607 8303 11633
rect 8329 11607 8386 11633
rect 8302 11606 8386 11607
rect 8302 11601 8330 11606
rect 8190 11159 8191 11185
rect 8217 11159 8218 11185
rect 8190 11153 8218 11159
rect 8246 11577 8274 11583
rect 8246 11551 8247 11577
rect 8273 11551 8274 11577
rect 8246 11466 8274 11551
rect 8134 11130 8162 11135
rect 8078 11102 8134 11130
rect 7854 11073 7882 11079
rect 7854 11047 7855 11073
rect 7881 11047 7882 11073
rect 7854 10906 7882 11047
rect 8022 10906 8050 10911
rect 7854 10878 8022 10906
rect 8022 10859 8050 10878
rect 7462 10431 7463 10457
rect 7489 10431 7490 10457
rect 7462 10425 7490 10431
rect 7518 10793 7658 10794
rect 7518 10767 7631 10793
rect 7657 10767 7658 10793
rect 7518 10766 7658 10767
rect 6062 9953 6090 10374
rect 6902 10402 6930 10407
rect 6902 10355 6930 10374
rect 6958 10402 6986 10407
rect 7070 10402 7098 10407
rect 6958 10401 7098 10402
rect 6958 10375 6959 10401
rect 6985 10375 7071 10401
rect 7097 10375 7098 10401
rect 6958 10374 7098 10375
rect 6958 10369 6986 10374
rect 7070 10369 7098 10374
rect 7350 10402 7378 10407
rect 7350 10401 7434 10402
rect 7350 10375 7351 10401
rect 7377 10375 7434 10401
rect 7350 10374 7434 10375
rect 7350 10369 7378 10374
rect 7238 10346 7266 10351
rect 7238 10299 7266 10318
rect 7350 10289 7378 10295
rect 7350 10263 7351 10289
rect 7377 10263 7378 10289
rect 7350 10178 7378 10263
rect 7126 10150 7378 10178
rect 7126 10065 7154 10150
rect 7126 10039 7127 10065
rect 7153 10039 7154 10065
rect 7126 10033 7154 10039
rect 6062 9927 6063 9953
rect 6089 9927 6090 9953
rect 6062 9921 6090 9927
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 966 9673 994 9679
rect 966 9647 967 9673
rect 993 9647 994 9673
rect 966 9450 994 9647
rect 2142 9618 2170 9623
rect 2142 9571 2170 9590
rect 6230 9618 6258 9623
rect 966 9417 994 9422
rect 6230 9169 6258 9590
rect 7294 9506 7322 9511
rect 6230 9143 6231 9169
rect 6257 9143 6258 9169
rect 6230 9137 6258 9143
rect 7014 9226 7042 9231
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 2142 8610 2170 8615
rect 2142 8441 2170 8582
rect 7014 8442 7042 9198
rect 7294 9225 7322 9478
rect 7406 9282 7434 10374
rect 7406 9249 7434 9254
rect 7518 10009 7546 10766
rect 7630 10761 7658 10766
rect 7966 10681 7994 10687
rect 7966 10655 7967 10681
rect 7993 10655 7994 10681
rect 7518 9983 7519 10009
rect 7545 9983 7546 10009
rect 7294 9199 7295 9225
rect 7321 9199 7322 9225
rect 7294 9193 7322 9199
rect 7518 9226 7546 9983
rect 7574 10345 7602 10351
rect 7574 10319 7575 10345
rect 7601 10319 7602 10345
rect 7574 9954 7602 10319
rect 7910 10346 7938 10351
rect 7910 10121 7938 10318
rect 7910 10095 7911 10121
rect 7937 10095 7938 10121
rect 7910 10089 7938 10095
rect 7630 9954 7658 9959
rect 7574 9926 7630 9954
rect 7630 9921 7658 9926
rect 7854 9674 7882 9679
rect 7798 9646 7854 9674
rect 7798 9617 7826 9646
rect 7854 9641 7882 9646
rect 7798 9591 7799 9617
rect 7825 9591 7826 9617
rect 7798 9585 7826 9591
rect 7966 9561 7994 10655
rect 8078 10065 8106 11102
rect 8134 11083 8162 11102
rect 8134 10906 8162 10911
rect 8246 10906 8274 11438
rect 8134 10905 8274 10906
rect 8134 10879 8135 10905
rect 8161 10879 8274 10905
rect 8134 10878 8274 10879
rect 8302 10906 8330 10911
rect 8358 10906 8386 11606
rect 8638 11633 8722 11634
rect 8638 11607 8695 11633
rect 8721 11607 8722 11633
rect 8638 11606 8722 11607
rect 8638 11186 8666 11606
rect 8694 11601 8722 11606
rect 8750 11466 8778 11471
rect 8778 11438 8946 11466
rect 8750 11419 8778 11438
rect 8638 11185 8778 11186
rect 8638 11159 8639 11185
rect 8665 11159 8778 11185
rect 8638 11158 8778 11159
rect 8638 11153 8666 11158
rect 8330 10878 8386 10906
rect 8694 11073 8722 11079
rect 8694 11047 8695 11073
rect 8721 11047 8722 11073
rect 8694 10906 8722 11047
rect 8134 10873 8162 10878
rect 8302 10873 8330 10878
rect 8302 10793 8330 10799
rect 8302 10767 8303 10793
rect 8329 10767 8330 10793
rect 8078 10039 8079 10065
rect 8105 10039 8106 10065
rect 8078 10033 8106 10039
rect 8246 10065 8274 10071
rect 8246 10039 8247 10065
rect 8273 10039 8274 10065
rect 8246 9730 8274 10039
rect 8302 10010 8330 10767
rect 8694 10793 8722 10878
rect 8694 10767 8695 10793
rect 8721 10767 8722 10793
rect 8694 10761 8722 10767
rect 8750 10794 8778 11158
rect 8918 11185 8946 11438
rect 8918 11159 8919 11185
rect 8945 11159 8946 11185
rect 8918 11153 8946 11159
rect 9086 11354 9114 11359
rect 8974 11130 9002 11135
rect 8974 11083 9002 11102
rect 8806 11074 8834 11079
rect 8806 11027 8834 11046
rect 9086 11073 9114 11326
rect 9086 11047 9087 11073
rect 9113 11047 9114 11073
rect 9086 10962 9114 11047
rect 9478 11074 9506 12335
rect 9590 12361 9618 12367
rect 9590 12335 9591 12361
rect 9617 12335 9618 12361
rect 9590 12250 9618 12335
rect 9590 12217 9618 12222
rect 9534 12026 9562 12031
rect 9646 12026 9674 13230
rect 10262 13257 10402 13258
rect 10262 13231 10263 13257
rect 10289 13231 10402 13257
rect 10262 13230 10402 13231
rect 10262 13225 10290 13230
rect 10318 13145 10346 13151
rect 10318 13119 10319 13145
rect 10345 13119 10346 13145
rect 9814 13034 9842 13039
rect 9814 12361 9842 13006
rect 10262 13034 10290 13039
rect 10262 12987 10290 13006
rect 10318 12922 10346 13119
rect 10262 12894 10346 12922
rect 10262 12698 10290 12894
rect 10318 12810 10346 12815
rect 10374 12810 10402 13230
rect 10318 12809 10402 12810
rect 10318 12783 10319 12809
rect 10345 12783 10402 12809
rect 10318 12782 10402 12783
rect 10318 12777 10346 12782
rect 10318 12698 10346 12703
rect 10262 12670 10318 12698
rect 10318 12665 10346 12670
rect 10542 12698 10570 12703
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12335 9815 12361
rect 9841 12335 9842 12361
rect 9814 12329 9842 12335
rect 10374 12362 10402 12367
rect 10374 12315 10402 12334
rect 9534 12025 9674 12026
rect 9534 11999 9535 12025
rect 9561 11999 9674 12025
rect 9534 11998 9674 11999
rect 9814 12250 9842 12255
rect 9534 11993 9562 11998
rect 9814 11970 9842 12222
rect 9814 11690 9842 11942
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9926 11690 9954 11695
rect 9814 11689 9954 11690
rect 9814 11663 9927 11689
rect 9953 11663 9954 11689
rect 9814 11662 9954 11663
rect 9926 11657 9954 11662
rect 10542 11689 10570 12670
rect 10542 11663 10543 11689
rect 10569 11663 10570 11689
rect 10542 11657 10570 11663
rect 10038 11577 10066 11583
rect 10038 11551 10039 11577
rect 10065 11551 10066 11577
rect 9870 11186 9898 11191
rect 9478 11041 9506 11046
rect 9646 11185 9898 11186
rect 9646 11159 9871 11185
rect 9897 11159 9898 11185
rect 9646 11158 9898 11159
rect 9086 10929 9114 10934
rect 9310 10906 9338 10911
rect 9254 10878 9310 10906
rect 8806 10794 8834 10799
rect 8750 10793 8834 10794
rect 8750 10767 8807 10793
rect 8833 10767 8834 10793
rect 8750 10766 8834 10767
rect 8806 10761 8834 10766
rect 8974 10682 9002 10687
rect 8974 10681 9114 10682
rect 8974 10655 8975 10681
rect 9001 10655 9114 10681
rect 8974 10654 9114 10655
rect 8974 10649 9002 10654
rect 8358 10010 8386 10015
rect 8302 10009 8386 10010
rect 8302 9983 8359 10009
rect 8385 9983 8386 10009
rect 8302 9982 8386 9983
rect 8358 9954 8386 9982
rect 9030 10010 9058 10015
rect 9030 9963 9058 9982
rect 8358 9921 8386 9926
rect 8246 9702 8386 9730
rect 8190 9674 8218 9679
rect 8190 9617 8218 9646
rect 8358 9674 8386 9702
rect 8190 9591 8191 9617
rect 8217 9591 8218 9617
rect 8190 9585 8218 9591
rect 8302 9618 8330 9623
rect 7966 9535 7967 9561
rect 7993 9535 7994 9561
rect 7854 9506 7882 9511
rect 7854 9459 7882 9478
rect 7686 9226 7714 9231
rect 7518 9198 7686 9226
rect 7686 9179 7714 9198
rect 7966 9170 7994 9535
rect 8078 9562 8106 9567
rect 8078 9515 8106 9534
rect 8302 9561 8330 9590
rect 8358 9617 8386 9646
rect 8358 9591 8359 9617
rect 8385 9591 8386 9617
rect 8358 9585 8386 9591
rect 8302 9535 8303 9561
rect 8329 9535 8330 9561
rect 8302 9529 8330 9535
rect 8750 9338 8778 9343
rect 8750 9291 8778 9310
rect 9030 9282 9058 9287
rect 8974 9254 9030 9282
rect 8918 9225 8946 9231
rect 8918 9199 8919 9225
rect 8945 9199 8946 9225
rect 7966 9137 7994 9142
rect 8862 9170 8890 9175
rect 8806 8890 8834 8895
rect 8134 8833 8162 8839
rect 8134 8807 8135 8833
rect 8161 8807 8162 8833
rect 7350 8722 7378 8727
rect 7294 8610 7322 8615
rect 2142 8415 2143 8441
rect 2169 8415 2170 8441
rect 2142 8409 2170 8415
rect 6790 8441 7042 8442
rect 6790 8415 7015 8441
rect 7041 8415 7042 8441
rect 6790 8414 7042 8415
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8073 994 8078
rect 6790 8049 6818 8414
rect 7014 8409 7042 8414
rect 7126 8498 7154 8503
rect 7126 8105 7154 8470
rect 7126 8079 7127 8105
rect 7153 8079 7154 8105
rect 7126 8073 7154 8079
rect 6790 8023 6791 8049
rect 6817 8023 6818 8049
rect 6790 8017 6818 8023
rect 7294 7769 7322 8582
rect 7350 8497 7378 8694
rect 7350 8471 7351 8497
rect 7377 8471 7378 8497
rect 7350 8465 7378 8471
rect 8134 8106 8162 8807
rect 8358 8833 8386 8839
rect 8358 8807 8359 8833
rect 8385 8807 8386 8833
rect 8358 8610 8386 8807
rect 8358 8577 8386 8582
rect 8414 8834 8442 8839
rect 8358 8442 8386 8447
rect 8190 8106 8218 8111
rect 8022 8105 8218 8106
rect 8022 8079 8191 8105
rect 8217 8079 8218 8105
rect 8022 8078 8218 8079
rect 7294 7743 7295 7769
rect 7321 7743 7322 7769
rect 7294 7658 7322 7743
rect 7630 7798 7994 7826
rect 7462 7714 7490 7719
rect 7462 7667 7490 7686
rect 7630 7713 7658 7798
rect 7630 7687 7631 7713
rect 7657 7687 7658 7713
rect 7630 7681 7658 7687
rect 7854 7714 7882 7719
rect 7294 7625 7322 7630
rect 7798 7658 7826 7663
rect 7798 7611 7826 7630
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 7742 2618 7770 2623
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 7406 1721 7434 1727
rect 7406 1695 7407 1721
rect 7433 1695 7434 1721
rect 4158 1666 4186 1671
rect 4046 1665 4186 1666
rect 4046 1639 4159 1665
rect 4185 1639 4186 1665
rect 4046 1638 4186 1639
rect 4046 400 4074 1638
rect 4158 1633 4186 1638
rect 7406 400 7434 1695
rect 7742 400 7770 2590
rect 7854 2561 7882 7686
rect 7854 2535 7855 2561
rect 7881 2535 7882 2561
rect 7854 2529 7882 2535
rect 7966 1777 7994 7798
rect 8022 7657 8050 8078
rect 8190 8073 8218 8078
rect 8302 8050 8330 8055
rect 8358 8050 8386 8414
rect 8414 8385 8442 8806
rect 8806 8833 8834 8862
rect 8806 8807 8807 8833
rect 8833 8807 8834 8833
rect 8806 8801 8834 8807
rect 8750 8498 8778 8503
rect 8750 8451 8778 8470
rect 8862 8497 8890 9142
rect 8918 8834 8946 9199
rect 8918 8801 8946 8806
rect 8918 8721 8946 8727
rect 8918 8695 8919 8721
rect 8945 8695 8946 8721
rect 8918 8666 8946 8695
rect 8918 8633 8946 8638
rect 8862 8471 8863 8497
rect 8889 8471 8890 8497
rect 8862 8465 8890 8471
rect 8974 8497 9002 9254
rect 9030 9249 9058 9254
rect 9086 8890 9114 10654
rect 9254 10066 9282 10878
rect 9310 10873 9338 10878
rect 9646 10849 9674 11158
rect 9870 11153 9898 11158
rect 9646 10823 9647 10849
rect 9673 10823 9674 10849
rect 9646 10817 9674 10823
rect 9814 11074 9842 11079
rect 9310 10794 9338 10799
rect 9310 10793 9394 10794
rect 9310 10767 9311 10793
rect 9337 10767 9394 10793
rect 9310 10766 9394 10767
rect 9310 10761 9338 10766
rect 9366 10345 9394 10766
rect 9366 10319 9367 10345
rect 9393 10319 9394 10345
rect 9254 10038 9338 10066
rect 9254 9954 9282 9959
rect 9254 9907 9282 9926
rect 9310 9618 9338 10038
rect 9310 9571 9338 9590
rect 9142 9562 9170 9567
rect 9142 9515 9170 9534
rect 9254 9506 9282 9511
rect 9254 9459 9282 9478
rect 9366 9394 9394 10319
rect 9814 10122 9842 11046
rect 9926 11074 9954 11093
rect 10038 11074 10066 11551
rect 10150 11186 10178 11191
rect 10598 11186 10626 11191
rect 10150 11185 10626 11186
rect 10150 11159 10151 11185
rect 10177 11159 10599 11185
rect 10625 11159 10626 11185
rect 10150 11158 10626 11159
rect 10150 11153 10178 11158
rect 10598 11153 10626 11158
rect 10654 11130 10682 15946
rect 11382 13258 11410 13263
rect 11382 13211 11410 13230
rect 11774 13258 11802 13263
rect 10822 13145 10850 13151
rect 10822 13119 10823 13145
rect 10849 13119 10850 13145
rect 10822 12642 10850 13119
rect 10934 13146 10962 13151
rect 11158 13146 11186 13151
rect 11270 13146 11298 13151
rect 10934 13145 11130 13146
rect 10934 13119 10935 13145
rect 10961 13119 11130 13145
rect 10934 13118 11130 13119
rect 10934 13113 10962 13118
rect 10822 12609 10850 12614
rect 10878 13089 10906 13095
rect 10878 13063 10879 13089
rect 10905 13063 10906 13089
rect 10710 12418 10738 12423
rect 10878 12418 10906 13063
rect 10710 12417 10906 12418
rect 10710 12391 10711 12417
rect 10737 12391 10906 12417
rect 10710 12390 10906 12391
rect 10934 12753 10962 12759
rect 10934 12727 10935 12753
rect 10961 12727 10962 12753
rect 10710 12385 10738 12390
rect 10934 12362 10962 12727
rect 10934 12329 10962 12334
rect 11046 12474 11074 12479
rect 10710 11578 10738 11583
rect 10710 11577 10794 11578
rect 10710 11551 10711 11577
rect 10737 11551 10794 11577
rect 10710 11550 10794 11551
rect 10710 11545 10738 11550
rect 10710 11130 10738 11135
rect 10654 11129 10738 11130
rect 10654 11103 10711 11129
rect 10737 11103 10738 11129
rect 10654 11102 10738 11103
rect 10038 11046 10122 11074
rect 9926 11041 9954 11046
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9814 10094 9898 10122
rect 9086 8833 9114 8862
rect 9254 9366 9394 9394
rect 9422 10009 9450 10015
rect 9422 9983 9423 10009
rect 9449 9983 9450 10009
rect 9422 9562 9450 9983
rect 9646 10010 9674 10015
rect 9646 9963 9674 9982
rect 9254 9226 9282 9366
rect 9366 9282 9394 9287
rect 9422 9282 9450 9534
rect 9534 9954 9562 9959
rect 9534 9561 9562 9926
rect 9758 9674 9786 9679
rect 9786 9646 9842 9674
rect 9758 9641 9786 9646
rect 9590 9618 9618 9623
rect 9618 9590 9674 9618
rect 9590 9585 9618 9590
rect 9534 9535 9535 9561
rect 9561 9535 9562 9561
rect 9534 9529 9562 9535
rect 9590 9506 9618 9511
rect 9366 9281 9450 9282
rect 9366 9255 9367 9281
rect 9393 9255 9450 9281
rect 9366 9254 9450 9255
rect 9478 9338 9506 9343
rect 9590 9338 9618 9478
rect 9646 9394 9674 9590
rect 9814 9561 9842 9646
rect 9870 9618 9898 10094
rect 10038 9674 10066 9679
rect 9982 9618 10010 9623
rect 9870 9617 10010 9618
rect 9870 9591 9983 9617
rect 10009 9591 10010 9617
rect 9870 9590 10010 9591
rect 9982 9585 10010 9590
rect 9814 9535 9815 9561
rect 9841 9535 9842 9561
rect 9646 9366 9786 9394
rect 9366 9249 9394 9254
rect 9086 8807 9087 8833
rect 9113 8807 9114 8833
rect 9086 8801 9114 8807
rect 9198 8834 9226 8839
rect 9198 8787 9226 8806
rect 8974 8471 8975 8497
rect 9001 8471 9002 8497
rect 8974 8465 9002 8471
rect 8638 8442 8666 8447
rect 8638 8395 8666 8414
rect 8414 8359 8415 8385
rect 8441 8359 8442 8385
rect 8414 8353 8442 8359
rect 8302 8049 8386 8050
rect 8302 8023 8303 8049
rect 8329 8023 8386 8049
rect 8302 8022 8386 8023
rect 8470 8050 8498 8055
rect 8302 8017 8330 8022
rect 8470 8003 8498 8022
rect 8414 7937 8442 7943
rect 8414 7911 8415 7937
rect 8441 7911 8442 7937
rect 8022 7631 8023 7657
rect 8049 7631 8050 7657
rect 8022 7625 8050 7631
rect 8134 7713 8162 7719
rect 8134 7687 8135 7713
rect 8161 7687 8162 7713
rect 7966 1751 7967 1777
rect 7993 1751 7994 1777
rect 7966 1745 7994 1751
rect 8134 1778 8162 7687
rect 8414 7658 8442 7911
rect 8414 7625 8442 7630
rect 9254 7657 9282 9198
rect 9478 9226 9506 9310
rect 9534 9310 9590 9338
rect 9534 9281 9562 9310
rect 9590 9305 9618 9310
rect 9534 9255 9535 9281
rect 9561 9255 9562 9281
rect 9534 9249 9562 9255
rect 9646 9282 9674 9287
rect 9646 9235 9674 9254
rect 9478 9193 9506 9198
rect 9702 9226 9730 9231
rect 9702 9179 9730 9198
rect 9310 9169 9338 9175
rect 9310 9143 9311 9169
rect 9337 9143 9338 9169
rect 9310 8834 9338 9143
rect 9310 8801 9338 8806
rect 9478 8834 9506 8839
rect 9478 8787 9506 8806
rect 9590 8833 9618 8839
rect 9590 8807 9591 8833
rect 9617 8807 9618 8833
rect 9590 8666 9618 8807
rect 9758 8833 9786 9366
rect 9814 9226 9842 9535
rect 9982 9506 10010 9511
rect 10038 9506 10066 9646
rect 9982 9505 10066 9506
rect 9982 9479 9983 9505
rect 10009 9479 10066 9505
rect 9982 9478 10066 9479
rect 9982 9473 10010 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10094 9394 10122 11046
rect 10710 10737 10738 11102
rect 10710 10711 10711 10737
rect 10737 10711 10738 10737
rect 10710 10705 10738 10711
rect 10766 11129 10794 11550
rect 10766 11103 10767 11129
rect 10793 11103 10794 11129
rect 10766 11074 10794 11103
rect 11046 11130 11074 12446
rect 11102 11970 11130 13118
rect 11158 13145 11298 13146
rect 11158 13119 11159 13145
rect 11185 13119 11271 13145
rect 11297 13119 11298 13145
rect 11158 13118 11298 13119
rect 11158 13113 11186 13118
rect 11270 13113 11298 13118
rect 11438 13145 11466 13151
rect 11438 13119 11439 13145
rect 11465 13119 11466 13145
rect 11270 12697 11298 12703
rect 11270 12671 11271 12697
rect 11297 12671 11298 12697
rect 11270 12026 11298 12671
rect 11438 12698 11466 13119
rect 11438 12665 11466 12670
rect 11774 12305 11802 13230
rect 12278 13258 12306 18999
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 12614 13454 12642 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12278 13225 12306 13230
rect 12334 13426 12642 13454
rect 12334 12810 12362 13426
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 11998 12809 12362 12810
rect 11998 12783 12335 12809
rect 12361 12783 12362 12809
rect 11998 12782 12362 12783
rect 11998 12473 12026 12782
rect 12334 12777 12362 12782
rect 13230 12698 13258 12703
rect 12166 12642 12194 12647
rect 11998 12447 11999 12473
rect 12025 12447 12026 12473
rect 11998 12441 12026 12447
rect 12054 12474 12082 12479
rect 12054 12417 12082 12446
rect 12054 12391 12055 12417
rect 12081 12391 12082 12417
rect 12054 12385 12082 12391
rect 11886 12362 11914 12367
rect 11774 12279 11775 12305
rect 11801 12279 11802 12305
rect 11774 12273 11802 12279
rect 11830 12361 11914 12362
rect 11830 12335 11887 12361
rect 11913 12335 11914 12361
rect 11830 12334 11914 12335
rect 11326 12026 11354 12031
rect 11830 12026 11858 12334
rect 11886 12329 11914 12334
rect 11270 12025 11354 12026
rect 11270 11999 11327 12025
rect 11353 11999 11354 12025
rect 11270 11998 11354 11999
rect 11326 11993 11354 11998
rect 11606 11998 11858 12026
rect 11130 11942 11298 11970
rect 11102 11923 11130 11942
rect 11270 11913 11298 11942
rect 11606 11969 11634 11998
rect 11606 11943 11607 11969
rect 11633 11943 11634 11969
rect 11606 11937 11634 11943
rect 11270 11887 11271 11913
rect 11297 11887 11298 11913
rect 11270 11881 11298 11887
rect 11382 11857 11410 11863
rect 11382 11831 11383 11857
rect 11409 11831 11410 11857
rect 11382 11354 11410 11831
rect 11382 11321 11410 11326
rect 12166 11857 12194 12614
rect 12502 12642 12530 12647
rect 12222 12306 12250 12311
rect 12222 12025 12250 12278
rect 12222 11999 12223 12025
rect 12249 11999 12250 12025
rect 12222 11993 12250 11999
rect 12502 11969 12530 12614
rect 13062 12642 13090 12647
rect 13062 12595 13090 12614
rect 13174 12641 13202 12647
rect 13174 12615 13175 12641
rect 13201 12615 13202 12641
rect 12502 11943 12503 11969
rect 12529 11943 12530 11969
rect 12502 11937 12530 11943
rect 12614 12362 12642 12367
rect 12614 11969 12642 12334
rect 13006 12306 13034 12311
rect 13006 12259 13034 12278
rect 13174 12306 13202 12615
rect 13174 12273 13202 12278
rect 12614 11943 12615 11969
rect 12641 11943 12642 11969
rect 12166 11831 12167 11857
rect 12193 11831 12194 11857
rect 11158 11130 11186 11135
rect 11046 11129 11186 11130
rect 11046 11103 11159 11129
rect 11185 11103 11186 11129
rect 11046 11102 11186 11103
rect 10990 11074 11018 11079
rect 10766 11073 11018 11074
rect 10766 11047 10991 11073
rect 11017 11047 11018 11073
rect 10766 11046 11018 11047
rect 10598 10346 10626 10351
rect 10626 10318 10682 10346
rect 10598 10313 10626 10318
rect 10206 9506 10234 9511
rect 10206 9459 10234 9478
rect 10374 9506 10402 9511
rect 10374 9459 10402 9478
rect 10094 9366 10346 9394
rect 10094 9338 10122 9366
rect 10094 9305 10122 9310
rect 9926 9282 9954 9287
rect 9870 9226 9898 9231
rect 9814 9225 9898 9226
rect 9814 9199 9871 9225
rect 9897 9199 9898 9225
rect 9814 9198 9898 9199
rect 9870 9114 9898 9198
rect 9870 9081 9898 9086
rect 9926 9002 9954 9254
rect 10318 9281 10346 9366
rect 10318 9255 10319 9281
rect 10345 9255 10346 9281
rect 10318 9249 10346 9255
rect 10598 9282 10626 9287
rect 9758 8807 9759 8833
rect 9785 8807 9786 8833
rect 9758 8778 9786 8807
rect 9758 8745 9786 8750
rect 9814 8974 9954 9002
rect 10094 9226 10122 9231
rect 9702 8722 9730 8727
rect 9702 8675 9730 8694
rect 9618 8638 9674 8666
rect 9590 8633 9618 8638
rect 9646 8554 9674 8638
rect 9702 8554 9730 8559
rect 9646 8553 9730 8554
rect 9646 8527 9703 8553
rect 9729 8527 9730 8553
rect 9646 8526 9730 8527
rect 9702 8442 9730 8526
rect 9814 8553 9842 8974
rect 9926 8834 9954 8839
rect 9926 8787 9954 8806
rect 10094 8777 10122 9198
rect 10150 9226 10178 9231
rect 10150 9225 10290 9226
rect 10150 9199 10151 9225
rect 10177 9199 10290 9225
rect 10150 9198 10290 9199
rect 10150 9193 10178 9198
rect 10094 8751 10095 8777
rect 10121 8751 10122 8777
rect 10094 8666 10122 8751
rect 10206 9114 10234 9119
rect 10206 8777 10234 9086
rect 10206 8751 10207 8777
rect 10233 8751 10234 8777
rect 10206 8745 10234 8751
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10094 8633 10122 8638
rect 10150 8721 10178 8727
rect 10150 8695 10151 8721
rect 10177 8695 10178 8721
rect 9918 8605 10050 8610
rect 9814 8527 9815 8553
rect 9841 8527 9842 8553
rect 9814 8521 9842 8527
rect 9982 8554 10010 8559
rect 10150 8554 10178 8695
rect 10262 8610 10290 9198
rect 10598 9225 10626 9254
rect 10598 9199 10599 9225
rect 10625 9199 10626 9225
rect 10598 9193 10626 9199
rect 10654 9170 10682 10318
rect 10766 9673 10794 11046
rect 10990 11041 11018 11046
rect 10822 10906 10850 10911
rect 10822 10457 10850 10878
rect 11158 10906 11186 11102
rect 11158 10873 11186 10878
rect 10990 10850 11018 10855
rect 10934 10793 10962 10799
rect 10934 10767 10935 10793
rect 10961 10767 10962 10793
rect 10934 10514 10962 10767
rect 10934 10481 10962 10486
rect 10822 10431 10823 10457
rect 10849 10431 10850 10457
rect 10822 10425 10850 10431
rect 10934 10402 10962 10407
rect 10990 10402 11018 10822
rect 12166 10850 12194 11831
rect 12278 11857 12306 11863
rect 12278 11831 12279 11857
rect 12305 11831 12306 11857
rect 12278 11690 12306 11831
rect 12278 11657 12306 11662
rect 12166 10817 12194 10822
rect 11270 10738 11298 10743
rect 12334 10738 12362 10743
rect 11270 10737 11690 10738
rect 11270 10711 11271 10737
rect 11297 10711 11690 10737
rect 11270 10710 11690 10711
rect 11270 10705 11298 10710
rect 10934 10401 11018 10402
rect 10934 10375 10935 10401
rect 10961 10375 11018 10401
rect 10934 10374 11018 10375
rect 11326 10402 11354 10407
rect 10934 10369 10962 10374
rect 11102 10290 11130 10295
rect 11102 10289 11298 10290
rect 11102 10263 11103 10289
rect 11129 10263 11298 10289
rect 11102 10262 11298 10263
rect 11102 10257 11130 10262
rect 11270 9898 11298 10262
rect 11326 10065 11354 10374
rect 11326 10039 11327 10065
rect 11353 10039 11354 10065
rect 11326 10033 11354 10039
rect 11270 9870 11578 9898
rect 10766 9647 10767 9673
rect 10793 9647 10794 9673
rect 10766 9641 10794 9647
rect 11550 9617 11578 9870
rect 11662 9673 11690 10710
rect 12278 10710 12334 10738
rect 11662 9647 11663 9673
rect 11689 9647 11690 9673
rect 11662 9641 11690 9647
rect 12054 9674 12082 9679
rect 11550 9591 11551 9617
rect 11577 9591 11578 9617
rect 11550 9585 11578 9591
rect 11774 9618 11802 9623
rect 11774 9571 11802 9590
rect 12054 9617 12082 9646
rect 12054 9591 12055 9617
rect 12081 9591 12082 9617
rect 12054 9585 12082 9591
rect 12110 9673 12138 9679
rect 12110 9647 12111 9673
rect 12137 9647 12138 9673
rect 12110 9618 12138 9647
rect 12110 9585 12138 9590
rect 10822 9562 10850 9567
rect 10990 9562 11018 9567
rect 10850 9561 11018 9562
rect 10850 9535 10991 9561
rect 11017 9535 11018 9561
rect 10850 9534 11018 9535
rect 10822 9515 10850 9534
rect 10990 9529 11018 9534
rect 11382 9562 11410 9567
rect 11382 9515 11410 9534
rect 11886 9561 11914 9567
rect 11886 9535 11887 9561
rect 11913 9535 11914 9561
rect 10710 9506 10738 9511
rect 10710 9459 10738 9478
rect 11046 9506 11074 9511
rect 10766 9338 10794 9343
rect 10766 9291 10794 9310
rect 11046 9337 11074 9478
rect 11158 9506 11186 9511
rect 11158 9459 11186 9478
rect 11214 9505 11242 9511
rect 11214 9479 11215 9505
rect 11241 9479 11242 9505
rect 11046 9311 11047 9337
rect 11073 9311 11074 9337
rect 11046 9305 11074 9311
rect 10822 9282 10850 9287
rect 10654 9142 10794 9170
rect 10654 8778 10682 8783
rect 10654 8731 10682 8750
rect 10262 8577 10290 8582
rect 10654 8610 10682 8615
rect 10206 8554 10234 8559
rect 9702 8409 9730 8414
rect 9926 8442 9954 8447
rect 9758 8385 9786 8391
rect 9758 8359 9759 8385
rect 9785 8359 9786 8385
rect 9254 7631 9255 7657
rect 9281 7631 9282 7657
rect 9254 7625 9282 7631
rect 9534 7938 9562 7943
rect 9534 6817 9562 7910
rect 9590 7714 9618 7719
rect 9758 7714 9786 8359
rect 9926 8105 9954 8414
rect 9982 8441 10010 8526
rect 9982 8415 9983 8441
rect 10009 8415 10010 8441
rect 9982 8409 10010 8415
rect 10094 8553 10234 8554
rect 10094 8527 10207 8553
rect 10233 8527 10234 8553
rect 10094 8526 10234 8527
rect 10094 8330 10122 8526
rect 10206 8521 10234 8526
rect 10318 8554 10346 8559
rect 10318 8507 10346 8526
rect 10150 8442 10178 8447
rect 10150 8395 10178 8414
rect 10094 8302 10178 8330
rect 9926 8079 9927 8105
rect 9953 8079 9954 8105
rect 9926 8073 9954 8079
rect 9814 8050 9842 8055
rect 9814 8003 9842 8022
rect 10150 8049 10178 8302
rect 10150 8023 10151 8049
rect 10177 8023 10178 8049
rect 10150 8017 10178 8023
rect 10598 8049 10626 8055
rect 10598 8023 10599 8049
rect 10625 8023 10626 8049
rect 10094 7994 10122 7999
rect 10038 7938 10066 7957
rect 10094 7947 10122 7966
rect 10598 7994 10626 8023
rect 10598 7961 10626 7966
rect 10038 7905 10066 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9590 7713 9786 7714
rect 9590 7687 9591 7713
rect 9617 7687 9786 7713
rect 9590 7686 9786 7687
rect 9590 7681 9618 7686
rect 10654 7601 10682 8582
rect 10766 8442 10794 9142
rect 10822 8833 10850 9254
rect 11214 9282 11242 9479
rect 11214 9249 11242 9254
rect 11326 9505 11354 9511
rect 11326 9479 11327 9505
rect 11353 9479 11354 9505
rect 10822 8807 10823 8833
rect 10849 8807 10850 8833
rect 10822 8801 10850 8807
rect 10878 9225 10906 9231
rect 10878 9199 10879 9225
rect 10905 9199 10906 9225
rect 10878 8834 10906 9199
rect 10878 8801 10906 8806
rect 11102 9170 11130 9175
rect 11326 9170 11354 9479
rect 11102 9169 11354 9170
rect 11102 9143 11103 9169
rect 11129 9143 11354 9169
rect 11102 9142 11354 9143
rect 11886 9338 11914 9535
rect 12278 9561 12306 10710
rect 12334 10691 12362 10710
rect 12614 10514 12642 11943
rect 13006 11914 13034 11919
rect 12726 11913 13034 11914
rect 12726 11887 13007 11913
rect 13033 11887 13034 11913
rect 12726 11886 13034 11887
rect 12614 10481 12642 10486
rect 12670 11690 12698 11695
rect 12670 10010 12698 11662
rect 12726 11689 12754 11886
rect 13006 11881 13034 11886
rect 12726 11663 12727 11689
rect 12753 11663 12754 11689
rect 12726 11657 12754 11663
rect 13230 11633 13258 12670
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 14070 12306 14098 12311
rect 14070 12259 14098 12278
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 13286 12026 13314 12031
rect 13286 11689 13314 11998
rect 14070 12026 14098 12031
rect 14070 11979 14098 11998
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 13286 11663 13287 11689
rect 13313 11663 13314 11689
rect 13286 11657 13314 11663
rect 13230 11607 13231 11633
rect 13257 11607 13258 11633
rect 13230 11601 13258 11607
rect 12782 11577 12810 11583
rect 12782 11551 12783 11577
rect 12809 11551 12810 11577
rect 12782 11354 12810 11551
rect 13006 11577 13034 11583
rect 13006 11551 13007 11577
rect 13033 11551 13034 11577
rect 13006 11466 13034 11551
rect 13286 11466 13314 11471
rect 13006 11465 13314 11466
rect 13006 11439 13287 11465
rect 13313 11439 13314 11465
rect 13006 11438 13314 11439
rect 13286 11433 13314 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 12782 11321 12810 11326
rect 13510 10906 13538 10911
rect 13062 10850 13090 10855
rect 13006 10849 13090 10850
rect 13006 10823 13063 10849
rect 13089 10823 13090 10849
rect 13006 10822 13090 10823
rect 12614 9982 12698 10010
rect 12726 10514 12754 10519
rect 12726 10345 12754 10486
rect 12726 10319 12727 10345
rect 12753 10319 12754 10345
rect 12726 10009 12754 10319
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12278 9535 12279 9561
rect 12305 9535 12306 9561
rect 12278 9529 12306 9535
rect 12446 9674 12474 9679
rect 12166 9506 12194 9511
rect 12166 9459 12194 9478
rect 11102 8610 11130 9142
rect 11774 8722 11802 8727
rect 11102 8577 11130 8582
rect 11606 8610 11634 8615
rect 10766 8049 10794 8414
rect 10766 8023 10767 8049
rect 10793 8023 10794 8049
rect 10766 8017 10794 8023
rect 10934 8498 10962 8503
rect 10934 8049 10962 8470
rect 11494 8498 11522 8503
rect 11494 8441 11522 8470
rect 11494 8415 11495 8441
rect 11521 8415 11522 8441
rect 11494 8409 11522 8415
rect 11606 8441 11634 8582
rect 11606 8415 11607 8441
rect 11633 8415 11634 8441
rect 11606 8409 11634 8415
rect 11774 8441 11802 8694
rect 11886 8498 11914 9310
rect 12054 8834 12082 8839
rect 12054 8787 12082 8806
rect 12334 8834 12362 8839
rect 12334 8787 12362 8806
rect 12446 8833 12474 9646
rect 12614 9337 12642 9982
rect 12726 9618 12754 9983
rect 13006 9674 13034 10822
rect 13062 10817 13090 10822
rect 13454 10849 13482 10855
rect 13454 10823 13455 10849
rect 13481 10823 13482 10849
rect 13118 10794 13146 10799
rect 13342 10794 13370 10799
rect 13118 10793 13370 10794
rect 13118 10767 13119 10793
rect 13145 10767 13343 10793
rect 13369 10767 13370 10793
rect 13118 10766 13370 10767
rect 13118 10761 13146 10766
rect 13342 10761 13370 10766
rect 13062 10681 13090 10687
rect 13062 10655 13063 10681
rect 13089 10655 13090 10681
rect 13062 10066 13090 10655
rect 13398 10514 13426 10519
rect 13118 10066 13146 10071
rect 13062 10065 13146 10066
rect 13062 10039 13119 10065
rect 13145 10039 13146 10065
rect 13062 10038 13146 10039
rect 13118 10033 13146 10038
rect 13006 9641 13034 9646
rect 12614 9311 12615 9337
rect 12641 9311 12642 9337
rect 12446 8807 12447 8833
rect 12473 8807 12474 8833
rect 12446 8801 12474 8807
rect 12558 8889 12586 8895
rect 12558 8863 12559 8889
rect 12585 8863 12586 8889
rect 12110 8722 12138 8727
rect 12110 8675 12138 8694
rect 12166 8721 12194 8727
rect 12166 8695 12167 8721
rect 12193 8695 12194 8721
rect 11886 8451 11914 8470
rect 11774 8415 11775 8441
rect 11801 8415 11802 8441
rect 11774 8409 11802 8415
rect 11998 8442 12026 8447
rect 11998 8395 12026 8414
rect 11662 8386 11690 8391
rect 11662 8339 11690 8358
rect 12054 8386 12082 8391
rect 11774 8050 11802 8055
rect 10934 8023 10935 8049
rect 10961 8023 10962 8049
rect 10934 8017 10962 8023
rect 11718 8022 11774 8050
rect 10654 7575 10655 7601
rect 10681 7575 10682 7601
rect 10654 7569 10682 7575
rect 10710 7937 10738 7943
rect 10710 7911 10711 7937
rect 10737 7911 10738 7937
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10598 6930 10626 6935
rect 10710 6930 10738 7911
rect 10990 7938 11018 7943
rect 10990 7769 11018 7910
rect 10990 7743 10991 7769
rect 11017 7743 11018 7769
rect 10990 7737 11018 7743
rect 10598 6929 10738 6930
rect 10598 6903 10599 6929
rect 10625 6903 10738 6929
rect 10598 6902 10738 6903
rect 10822 7713 10850 7719
rect 10822 7687 10823 7713
rect 10849 7687 10850 7713
rect 10598 6897 10626 6902
rect 9534 6791 9535 6817
rect 9561 6791 9562 6817
rect 9534 6706 9562 6791
rect 9534 6673 9562 6678
rect 10206 6706 10234 6711
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 8358 2618 8386 2623
rect 8358 2571 8386 2590
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10206 2169 10234 6678
rect 10206 2143 10207 2169
rect 10233 2143 10234 2169
rect 10206 2137 10234 2143
rect 10094 2058 10122 2063
rect 8470 1778 8498 1783
rect 8134 1777 8498 1778
rect 8134 1751 8471 1777
rect 8497 1751 8498 1777
rect 8134 1750 8498 1751
rect 8470 1745 8498 1750
rect 8078 1722 8106 1727
rect 8078 400 8106 1694
rect 9254 1722 9282 1727
rect 9254 1675 9282 1694
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10094 400 10122 2030
rect 10710 2058 10738 2063
rect 10710 2011 10738 2030
rect 10766 1834 10794 1839
rect 10766 400 10794 1806
rect 10822 1777 10850 7687
rect 10934 7602 10962 7607
rect 10934 6873 10962 7574
rect 11718 7602 11746 8022
rect 11774 8003 11802 8022
rect 11718 7265 11746 7574
rect 12054 7321 12082 8358
rect 12110 8385 12138 8391
rect 12110 8359 12111 8385
rect 12137 8359 12138 8385
rect 12110 8105 12138 8359
rect 12110 8079 12111 8105
rect 12137 8079 12138 8105
rect 12110 8073 12138 8079
rect 12166 7770 12194 8695
rect 12222 8498 12250 8503
rect 12222 8441 12250 8470
rect 12558 8498 12586 8863
rect 12614 8834 12642 9311
rect 12614 8787 12642 8806
rect 12670 9617 12754 9618
rect 12670 9591 12727 9617
rect 12753 9591 12754 9617
rect 12670 9590 12754 9591
rect 12558 8465 12586 8470
rect 12222 8415 12223 8441
rect 12249 8415 12250 8441
rect 12222 8409 12250 8415
rect 12670 8050 12698 9590
rect 12726 9585 12754 9590
rect 13118 9562 13146 9567
rect 13118 9561 13258 9562
rect 13118 9535 13119 9561
rect 13145 9535 13258 9561
rect 13118 9534 13258 9535
rect 13118 9529 13146 9534
rect 12726 9506 12754 9511
rect 12726 9225 12754 9478
rect 13230 9337 13258 9534
rect 13230 9311 13231 9337
rect 13257 9311 13258 9337
rect 13230 9305 13258 9311
rect 12726 9199 12727 9225
rect 12753 9199 12754 9225
rect 12726 9193 12754 9199
rect 13342 9281 13370 9287
rect 13342 9255 13343 9281
rect 13369 9255 13370 9281
rect 12726 8722 12754 8727
rect 12726 8675 12754 8694
rect 13118 8722 13146 8727
rect 13118 8553 13146 8694
rect 13342 8610 13370 9255
rect 13398 9281 13426 10486
rect 13454 10122 13482 10823
rect 13510 10849 13538 10878
rect 13510 10823 13511 10849
rect 13537 10823 13538 10849
rect 13510 10817 13538 10823
rect 14126 10906 14154 10911
rect 14126 10401 14154 10878
rect 18942 10793 18970 10799
rect 18942 10767 18943 10793
rect 18969 10767 18970 10793
rect 18830 10682 18858 10687
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 14182 10514 14210 10519
rect 14182 10467 14210 10486
rect 14126 10375 14127 10401
rect 14153 10375 14154 10401
rect 14126 10369 14154 10375
rect 18830 10401 18858 10654
rect 18830 10375 18831 10401
rect 18857 10375 18858 10401
rect 18830 10369 18858 10375
rect 14182 10290 14210 10295
rect 14182 10289 14266 10290
rect 14182 10263 14183 10289
rect 14209 10263 14266 10289
rect 14182 10262 14266 10263
rect 14182 10257 14210 10262
rect 13454 10089 13482 10094
rect 14182 10122 14210 10127
rect 14182 9953 14210 10094
rect 14182 9927 14183 9953
rect 14209 9927 14210 9953
rect 14182 9921 14210 9927
rect 13398 9255 13399 9281
rect 13425 9255 13426 9281
rect 13398 9249 13426 9255
rect 14238 9505 14266 10262
rect 18942 10122 18970 10767
rect 19950 10737 19978 10743
rect 19950 10711 19951 10737
rect 19977 10711 19978 10737
rect 19950 10458 19978 10711
rect 19950 10425 19978 10430
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 18942 10089 18970 10094
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 18830 10010 18858 10015
rect 18774 10009 18858 10010
rect 18774 9983 18831 10009
rect 18857 9983 18858 10009
rect 18774 9982 18858 9983
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 14238 9479 14239 9505
rect 14265 9479 14266 9505
rect 14238 9282 14266 9479
rect 14630 9617 14658 9623
rect 14630 9591 14631 9617
rect 14657 9591 14658 9617
rect 14350 9282 14378 9287
rect 14238 9254 14350 9282
rect 14350 9225 14378 9254
rect 14350 9199 14351 9225
rect 14377 9199 14378 9225
rect 14350 9193 14378 9199
rect 14462 9281 14490 9287
rect 14462 9255 14463 9281
rect 14489 9255 14490 9281
rect 14462 9226 14490 9255
rect 14630 9282 14658 9591
rect 14742 9506 14770 9511
rect 14742 9459 14770 9478
rect 14630 9249 14658 9254
rect 14462 9193 14490 9198
rect 18774 9226 18802 9982
rect 18830 9977 18858 9982
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 18830 9617 18858 9623
rect 18830 9591 18831 9617
rect 18857 9591 18858 9617
rect 18830 9338 18858 9591
rect 18830 9305 18858 9310
rect 18942 9506 18970 9511
rect 18774 9193 18802 9198
rect 18942 9225 18970 9478
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 18942 9199 18943 9225
rect 18969 9199 18970 9225
rect 18942 9193 18970 9199
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 13342 8577 13370 8582
rect 18942 8833 18970 8839
rect 18942 8807 18943 8833
rect 18969 8807 18970 8833
rect 13118 8527 13119 8553
rect 13145 8527 13146 8553
rect 13118 8442 13146 8527
rect 13286 8497 13314 8503
rect 13286 8471 13287 8497
rect 13313 8471 13314 8497
rect 13146 8414 13202 8442
rect 13118 8409 13146 8414
rect 13174 8105 13202 8414
rect 13286 8386 13314 8471
rect 13286 8353 13314 8358
rect 18830 8441 18858 8447
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 18830 8386 18858 8415
rect 18942 8442 18970 8807
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 18942 8409 18970 8414
rect 20006 8442 20034 8447
rect 18830 8353 18858 8358
rect 20006 8385 20034 8414
rect 20006 8359 20007 8385
rect 20033 8359 20034 8385
rect 20006 8353 20034 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 13174 8079 13175 8105
rect 13201 8079 13202 8105
rect 13174 8073 13202 8079
rect 20006 8106 20034 8111
rect 20006 8059 20034 8078
rect 12670 8017 12698 8022
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 12166 7737 12194 7742
rect 12782 7770 12810 7775
rect 12054 7295 12055 7321
rect 12081 7295 12082 7321
rect 12054 7289 12082 7295
rect 12782 7322 12810 7742
rect 12950 7714 12978 7719
rect 12950 7667 12978 7686
rect 18830 7714 18858 8023
rect 18830 7681 18858 7686
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13118 7322 13146 7327
rect 12782 7321 13146 7322
rect 12782 7295 13119 7321
rect 13145 7295 13146 7321
rect 12782 7294 13146 7295
rect 11718 7239 11719 7265
rect 11745 7239 11746 7265
rect 11718 7233 11746 7239
rect 10934 6847 10935 6873
rect 10961 6847 10962 6873
rect 10934 6841 10962 6847
rect 12782 4214 12810 7294
rect 13118 7289 13146 7294
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 12614 4186 12810 4214
rect 11214 1834 11242 1839
rect 11214 1787 11242 1806
rect 12446 1834 12474 1839
rect 10822 1751 10823 1777
rect 10849 1751 10850 1777
rect 10822 1745 10850 1751
rect 12446 400 12474 1806
rect 12614 1777 12642 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 13062 1834 13090 1839
rect 13062 1787 13090 1806
rect 12614 1751 12615 1777
rect 12641 1751 12642 1777
rect 12614 1745 12642 1751
rect 15246 1666 15274 1671
rect 15134 1665 15274 1666
rect 15134 1639 15247 1665
rect 15273 1639 15274 1665
rect 15134 1638 15274 1639
rect 15134 400 15162 1638
rect 15246 1633 15274 1638
rect 4032 0 4088 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 10080 0 10136 400
rect 10752 0 10808 400
rect 12432 0 12488 400
rect 15120 0 15176 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 10766 19110 10794 19138
rect 11214 19137 11242 19138
rect 11214 19111 11215 19137
rect 11215 19111 11241 19137
rect 11241 19111 11242 19137
rect 11214 19110 11242 19111
rect 11774 19110 11802 19138
rect 10430 18718 10458 18746
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 11046 18745 11074 18746
rect 11046 18719 11047 18745
rect 11047 18719 11073 18745
rect 11073 18719 11074 18745
rect 11046 18718 11074 18719
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 12110 18718 12138 18746
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9086 13006 9114 13034
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2086 12782 2114 12810
rect 966 10430 994 10458
rect 7238 12614 7266 12642
rect 6902 12390 6930 12418
rect 8078 12641 8106 12642
rect 8078 12615 8079 12641
rect 8079 12615 8105 12641
rect 8105 12615 8106 12641
rect 8078 12614 8106 12615
rect 8190 12641 8218 12642
rect 8190 12615 8191 12641
rect 8191 12615 8217 12641
rect 8217 12615 8218 12641
rect 8190 12614 8218 12615
rect 7630 12390 7658 12418
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6174 11158 6202 11186
rect 2142 10793 2170 10794
rect 2142 10767 2143 10793
rect 2143 10767 2169 10793
rect 2169 10767 2170 10793
rect 2142 10766 2170 10767
rect 6062 10766 6090 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2086 9926 2114 9954
rect 7462 11185 7490 11186
rect 7462 11159 7463 11185
rect 7463 11159 7489 11185
rect 7489 11159 7490 11185
rect 7462 11158 7490 11159
rect 7406 11102 7434 11130
rect 7462 10934 7490 10962
rect 8134 12390 8162 12418
rect 8862 12390 8890 12418
rect 8358 12334 8386 12362
rect 8302 11718 8330 11746
rect 7686 11185 7714 11186
rect 7686 11159 7687 11185
rect 7687 11159 7713 11185
rect 7713 11159 7714 11185
rect 7686 11158 7714 11159
rect 8806 12361 8834 12362
rect 8806 12335 8807 12361
rect 8807 12335 8833 12361
rect 8833 12335 8834 12361
rect 8806 12334 8834 12335
rect 9534 13033 9562 13034
rect 9534 13007 9535 13033
rect 9535 13007 9561 13033
rect 9561 13007 9562 13033
rect 9534 13006 9562 13007
rect 9590 12446 9618 12474
rect 8918 12222 8946 12250
rect 8694 11718 8722 11746
rect 8246 11438 8274 11466
rect 8134 11129 8162 11130
rect 8134 11103 8135 11129
rect 8135 11103 8161 11129
rect 8161 11103 8162 11129
rect 8134 11102 8162 11103
rect 8022 10905 8050 10906
rect 8022 10879 8023 10905
rect 8023 10879 8049 10905
rect 8049 10879 8050 10905
rect 8022 10878 8050 10879
rect 6062 10374 6090 10402
rect 6902 10401 6930 10402
rect 6902 10375 6903 10401
rect 6903 10375 6929 10401
rect 6929 10375 6930 10401
rect 6902 10374 6930 10375
rect 7238 10345 7266 10346
rect 7238 10319 7239 10345
rect 7239 10319 7265 10345
rect 7265 10319 7266 10345
rect 7238 10318 7266 10319
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 2142 9617 2170 9618
rect 2142 9591 2143 9617
rect 2143 9591 2169 9617
rect 2169 9591 2170 9617
rect 2142 9590 2170 9591
rect 6230 9590 6258 9618
rect 966 9422 994 9450
rect 7294 9478 7322 9506
rect 7014 9198 7042 9226
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2142 8582 2170 8610
rect 7406 9254 7434 9282
rect 7910 10318 7938 10346
rect 7630 9926 7658 9954
rect 7854 9646 7882 9674
rect 8750 11465 8778 11466
rect 8750 11439 8751 11465
rect 8751 11439 8777 11465
rect 8777 11439 8778 11465
rect 8750 11438 8778 11439
rect 8302 10878 8330 10906
rect 8694 10878 8722 10906
rect 9086 11326 9114 11354
rect 8974 11129 9002 11130
rect 8974 11103 8975 11129
rect 8975 11103 9001 11129
rect 9001 11103 9002 11129
rect 8974 11102 9002 11103
rect 8806 11073 8834 11074
rect 8806 11047 8807 11073
rect 8807 11047 8833 11073
rect 8833 11047 8834 11073
rect 8806 11046 8834 11047
rect 9590 12222 9618 12250
rect 9814 13006 9842 13034
rect 10262 13033 10290 13034
rect 10262 13007 10263 13033
rect 10263 13007 10289 13033
rect 10289 13007 10290 13033
rect 10262 13006 10290 13007
rect 10318 12670 10346 12698
rect 10542 12670 10570 12698
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10374 12361 10402 12362
rect 10374 12335 10375 12361
rect 10375 12335 10401 12361
rect 10401 12335 10402 12361
rect 10374 12334 10402 12335
rect 9814 12222 9842 12250
rect 9814 11942 9842 11970
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9478 11046 9506 11074
rect 9086 10934 9114 10962
rect 9310 10878 9338 10906
rect 9030 10009 9058 10010
rect 9030 9983 9031 10009
rect 9031 9983 9057 10009
rect 9057 9983 9058 10009
rect 9030 9982 9058 9983
rect 8358 9926 8386 9954
rect 8190 9646 8218 9674
rect 8358 9646 8386 9674
rect 8302 9590 8330 9618
rect 7854 9505 7882 9506
rect 7854 9479 7855 9505
rect 7855 9479 7881 9505
rect 7881 9479 7882 9505
rect 7854 9478 7882 9479
rect 7686 9225 7714 9226
rect 7686 9199 7687 9225
rect 7687 9199 7713 9225
rect 7713 9199 7714 9225
rect 7686 9198 7714 9199
rect 8078 9561 8106 9562
rect 8078 9535 8079 9561
rect 8079 9535 8105 9561
rect 8105 9535 8106 9561
rect 8078 9534 8106 9535
rect 8750 9337 8778 9338
rect 8750 9311 8751 9337
rect 8751 9311 8777 9337
rect 8777 9311 8778 9337
rect 8750 9310 8778 9311
rect 9030 9254 9058 9282
rect 7966 9142 7994 9170
rect 8862 9142 8890 9170
rect 8806 8862 8834 8890
rect 7350 8694 7378 8722
rect 7294 8582 7322 8610
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 966 8078 994 8106
rect 7126 8470 7154 8498
rect 8358 8582 8386 8610
rect 8414 8806 8442 8834
rect 8358 8414 8386 8442
rect 7462 7713 7490 7714
rect 7462 7687 7463 7713
rect 7463 7687 7489 7713
rect 7489 7687 7490 7713
rect 7462 7686 7490 7687
rect 7854 7686 7882 7714
rect 7294 7630 7322 7658
rect 7798 7657 7826 7658
rect 7798 7631 7799 7657
rect 7799 7631 7825 7657
rect 7825 7631 7826 7657
rect 7798 7630 7826 7631
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 7742 2590 7770 2618
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 8750 8497 8778 8498
rect 8750 8471 8751 8497
rect 8751 8471 8777 8497
rect 8777 8471 8778 8497
rect 8750 8470 8778 8471
rect 8918 8806 8946 8834
rect 8918 8638 8946 8666
rect 9814 11073 9842 11074
rect 9814 11047 9815 11073
rect 9815 11047 9841 11073
rect 9841 11047 9842 11073
rect 9814 11046 9842 11047
rect 9254 9953 9282 9954
rect 9254 9927 9255 9953
rect 9255 9927 9281 9953
rect 9281 9927 9282 9953
rect 9254 9926 9282 9927
rect 9310 9617 9338 9618
rect 9310 9591 9311 9617
rect 9311 9591 9337 9617
rect 9337 9591 9338 9617
rect 9310 9590 9338 9591
rect 9142 9561 9170 9562
rect 9142 9535 9143 9561
rect 9143 9535 9169 9561
rect 9169 9535 9170 9561
rect 9142 9534 9170 9535
rect 9254 9505 9282 9506
rect 9254 9479 9255 9505
rect 9255 9479 9281 9505
rect 9281 9479 9282 9505
rect 9254 9478 9282 9479
rect 9926 11073 9954 11074
rect 9926 11047 9927 11073
rect 9927 11047 9953 11073
rect 9953 11047 9954 11073
rect 9926 11046 9954 11047
rect 11382 13257 11410 13258
rect 11382 13231 11383 13257
rect 11383 13231 11409 13257
rect 11409 13231 11410 13257
rect 11382 13230 11410 13231
rect 11774 13230 11802 13258
rect 10822 12614 10850 12642
rect 10934 12334 10962 12362
rect 11046 12446 11074 12474
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9086 8862 9114 8890
rect 9646 10009 9674 10010
rect 9646 9983 9647 10009
rect 9647 9983 9673 10009
rect 9673 9983 9674 10009
rect 9646 9982 9674 9983
rect 9422 9534 9450 9562
rect 9534 9926 9562 9954
rect 9758 9646 9786 9674
rect 9590 9590 9618 9618
rect 9590 9478 9618 9506
rect 10038 9646 10066 9674
rect 9478 9310 9506 9338
rect 9254 9198 9282 9226
rect 9198 8833 9226 8834
rect 9198 8807 9199 8833
rect 9199 8807 9225 8833
rect 9225 8807 9226 8833
rect 9198 8806 9226 8807
rect 8638 8441 8666 8442
rect 8638 8415 8639 8441
rect 8639 8415 8665 8441
rect 8665 8415 8666 8441
rect 8638 8414 8666 8415
rect 8470 8049 8498 8050
rect 8470 8023 8471 8049
rect 8471 8023 8497 8049
rect 8497 8023 8498 8049
rect 8470 8022 8498 8023
rect 8414 7630 8442 7658
rect 9590 9310 9618 9338
rect 9646 9281 9674 9282
rect 9646 9255 9647 9281
rect 9647 9255 9673 9281
rect 9673 9255 9674 9281
rect 9646 9254 9674 9255
rect 9478 9198 9506 9226
rect 9702 9225 9730 9226
rect 9702 9199 9703 9225
rect 9703 9199 9729 9225
rect 9729 9199 9730 9225
rect 9702 9198 9730 9199
rect 9310 8806 9338 8834
rect 9478 8833 9506 8834
rect 9478 8807 9479 8833
rect 9479 8807 9505 8833
rect 9505 8807 9506 8833
rect 9478 8806 9506 8807
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 11438 12670 11466 12698
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12278 13230 12306 13258
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 13230 12697 13258 12698
rect 13230 12671 13231 12697
rect 13231 12671 13257 12697
rect 13257 12671 13258 12697
rect 13230 12670 13258 12671
rect 12166 12614 12194 12642
rect 12054 12446 12082 12474
rect 11102 11942 11130 11970
rect 11382 11326 11410 11354
rect 12502 12614 12530 12642
rect 12222 12278 12250 12306
rect 13062 12641 13090 12642
rect 13062 12615 13063 12641
rect 13063 12615 13089 12641
rect 13089 12615 13090 12641
rect 13062 12614 13090 12615
rect 12614 12361 12642 12362
rect 12614 12335 12615 12361
rect 12615 12335 12641 12361
rect 12641 12335 12642 12361
rect 12614 12334 12642 12335
rect 13006 12305 13034 12306
rect 13006 12279 13007 12305
rect 13007 12279 13033 12305
rect 13033 12279 13034 12305
rect 13006 12278 13034 12279
rect 13174 12278 13202 12306
rect 10598 10318 10626 10346
rect 10206 9505 10234 9506
rect 10206 9479 10207 9505
rect 10207 9479 10233 9505
rect 10233 9479 10234 9505
rect 10206 9478 10234 9479
rect 10374 9505 10402 9506
rect 10374 9479 10375 9505
rect 10375 9479 10401 9505
rect 10401 9479 10402 9505
rect 10374 9478 10402 9479
rect 10094 9310 10122 9338
rect 9926 9254 9954 9282
rect 9870 9086 9898 9114
rect 10598 9254 10626 9282
rect 9758 8750 9786 8778
rect 10094 9198 10122 9226
rect 9702 8721 9730 8722
rect 9702 8695 9703 8721
rect 9703 8695 9729 8721
rect 9729 8695 9730 8721
rect 9702 8694 9730 8695
rect 9590 8638 9618 8666
rect 9926 8833 9954 8834
rect 9926 8807 9927 8833
rect 9927 8807 9953 8833
rect 9953 8807 9954 8833
rect 9926 8806 9954 8807
rect 10206 9086 10234 9114
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10094 8638 10122 8666
rect 10022 8610 10050 8611
rect 10822 10878 10850 10906
rect 11158 10878 11186 10906
rect 10990 10822 11018 10850
rect 10934 10486 10962 10514
rect 12278 11662 12306 11690
rect 12166 10822 12194 10850
rect 11326 10401 11354 10402
rect 11326 10375 11327 10401
rect 11327 10375 11353 10401
rect 11353 10375 11354 10401
rect 11326 10374 11354 10375
rect 12334 10737 12362 10738
rect 12334 10711 12335 10737
rect 12335 10711 12361 10737
rect 12361 10711 12362 10737
rect 12334 10710 12362 10711
rect 12054 9646 12082 9674
rect 11774 9617 11802 9618
rect 11774 9591 11775 9617
rect 11775 9591 11801 9617
rect 11801 9591 11802 9617
rect 11774 9590 11802 9591
rect 12110 9590 12138 9618
rect 10822 9561 10850 9562
rect 10822 9535 10823 9561
rect 10823 9535 10849 9561
rect 10849 9535 10850 9561
rect 10822 9534 10850 9535
rect 11382 9561 11410 9562
rect 11382 9535 11383 9561
rect 11383 9535 11409 9561
rect 11409 9535 11410 9561
rect 11382 9534 11410 9535
rect 10710 9505 10738 9506
rect 10710 9479 10711 9505
rect 10711 9479 10737 9505
rect 10737 9479 10738 9505
rect 10710 9478 10738 9479
rect 11046 9505 11074 9506
rect 11046 9479 11047 9505
rect 11047 9479 11073 9505
rect 11073 9479 11074 9505
rect 11046 9478 11074 9479
rect 10766 9337 10794 9338
rect 10766 9311 10767 9337
rect 10767 9311 10793 9337
rect 10793 9311 10794 9337
rect 10766 9310 10794 9311
rect 11158 9505 11186 9506
rect 11158 9479 11159 9505
rect 11159 9479 11185 9505
rect 11185 9479 11186 9505
rect 11158 9478 11186 9479
rect 10822 9254 10850 9282
rect 10654 8777 10682 8778
rect 10654 8751 10655 8777
rect 10655 8751 10681 8777
rect 10681 8751 10682 8777
rect 10654 8750 10682 8751
rect 10262 8582 10290 8610
rect 10654 8582 10682 8610
rect 9982 8526 10010 8554
rect 9702 8414 9730 8442
rect 9926 8414 9954 8442
rect 9534 7910 9562 7938
rect 10318 8553 10346 8554
rect 10318 8527 10319 8553
rect 10319 8527 10345 8553
rect 10345 8527 10346 8553
rect 10318 8526 10346 8527
rect 10150 8441 10178 8442
rect 10150 8415 10151 8441
rect 10151 8415 10177 8441
rect 10177 8415 10178 8441
rect 10150 8414 10178 8415
rect 9814 8049 9842 8050
rect 9814 8023 9815 8049
rect 9815 8023 9841 8049
rect 9841 8023 9842 8049
rect 9814 8022 9842 8023
rect 10094 7993 10122 7994
rect 10094 7967 10095 7993
rect 10095 7967 10121 7993
rect 10121 7967 10122 7993
rect 10094 7966 10122 7967
rect 10598 7966 10626 7994
rect 10038 7937 10066 7938
rect 10038 7911 10039 7937
rect 10039 7911 10065 7937
rect 10065 7911 10066 7937
rect 10038 7910 10066 7911
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 11214 9254 11242 9282
rect 10878 8806 10906 8834
rect 12614 10486 12642 10514
rect 12670 11689 12698 11690
rect 12670 11663 12671 11689
rect 12671 11663 12697 11689
rect 12697 11663 12698 11689
rect 12670 11662 12698 11663
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 14070 12305 14098 12306
rect 14070 12279 14071 12305
rect 14071 12279 14097 12305
rect 14097 12279 14098 12305
rect 14070 12278 14098 12279
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 13286 11998 13314 12026
rect 14070 12025 14098 12026
rect 14070 11999 14071 12025
rect 14071 11999 14097 12025
rect 14097 11999 14098 12025
rect 14070 11998 14098 11999
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 20006 11774 20034 11802
rect 12782 11326 12810 11354
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 13510 10878 13538 10906
rect 12726 10486 12754 10514
rect 12446 9646 12474 9674
rect 12166 9505 12194 9506
rect 12166 9479 12167 9505
rect 12167 9479 12193 9505
rect 12193 9479 12194 9505
rect 12166 9478 12194 9479
rect 11886 9310 11914 9338
rect 11774 8694 11802 8722
rect 11102 8582 11130 8610
rect 11606 8582 11634 8610
rect 10766 8414 10794 8442
rect 10934 8470 10962 8498
rect 11494 8470 11522 8498
rect 12054 8833 12082 8834
rect 12054 8807 12055 8833
rect 12055 8807 12081 8833
rect 12081 8807 12082 8833
rect 12054 8806 12082 8807
rect 12334 8833 12362 8834
rect 12334 8807 12335 8833
rect 12335 8807 12361 8833
rect 12361 8807 12362 8833
rect 12334 8806 12362 8807
rect 13398 10486 13426 10514
rect 13006 9646 13034 9674
rect 12110 8721 12138 8722
rect 12110 8695 12111 8721
rect 12111 8695 12137 8721
rect 12137 8695 12138 8721
rect 12110 8694 12138 8695
rect 11886 8497 11914 8498
rect 11886 8471 11887 8497
rect 11887 8471 11913 8497
rect 11913 8471 11914 8497
rect 11886 8470 11914 8471
rect 11998 8441 12026 8442
rect 11998 8415 11999 8441
rect 11999 8415 12025 8441
rect 12025 8415 12026 8441
rect 11998 8414 12026 8415
rect 11662 8385 11690 8386
rect 11662 8359 11663 8385
rect 11663 8359 11689 8385
rect 11689 8359 11690 8385
rect 11662 8358 11690 8359
rect 12054 8358 12082 8386
rect 11774 8049 11802 8050
rect 11774 8023 11775 8049
rect 11775 8023 11801 8049
rect 11801 8023 11802 8049
rect 11774 8022 11802 8023
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10990 7910 11018 7938
rect 9534 6678 9562 6706
rect 10206 6678 10234 6706
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 8358 2617 8386 2618
rect 8358 2591 8359 2617
rect 8359 2591 8385 2617
rect 8385 2591 8386 2617
rect 8358 2590 8386 2591
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 10094 2030 10122 2058
rect 8078 1694 8106 1722
rect 9254 1721 9282 1722
rect 9254 1695 9255 1721
rect 9255 1695 9281 1721
rect 9281 1695 9282 1721
rect 9254 1694 9282 1695
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 10710 2057 10738 2058
rect 10710 2031 10711 2057
rect 10711 2031 10737 2057
rect 10737 2031 10738 2057
rect 10710 2030 10738 2031
rect 10766 1806 10794 1834
rect 10934 7574 10962 7602
rect 11718 7574 11746 7602
rect 12222 8470 12250 8498
rect 12614 8833 12642 8834
rect 12614 8807 12615 8833
rect 12615 8807 12641 8833
rect 12641 8807 12642 8833
rect 12614 8806 12642 8807
rect 12558 8470 12586 8498
rect 12726 9478 12754 9506
rect 12726 8721 12754 8722
rect 12726 8695 12727 8721
rect 12727 8695 12753 8721
rect 12753 8695 12754 8721
rect 12726 8694 12754 8695
rect 13118 8694 13146 8722
rect 14126 10878 14154 10906
rect 18830 10654 18858 10682
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 14182 10513 14210 10514
rect 14182 10487 14183 10513
rect 14183 10487 14209 10513
rect 14209 10487 14210 10513
rect 14182 10486 14210 10487
rect 13454 10094 13482 10122
rect 14182 10094 14210 10122
rect 19950 10430 19978 10458
rect 18942 10094 18970 10122
rect 20006 10094 20034 10122
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14350 9254 14378 9282
rect 14742 9505 14770 9506
rect 14742 9479 14743 9505
rect 14743 9479 14769 9505
rect 14769 9479 14770 9505
rect 14742 9478 14770 9479
rect 14630 9254 14658 9282
rect 14462 9198 14490 9226
rect 20006 9758 20034 9786
rect 18830 9310 18858 9338
rect 18942 9478 18970 9506
rect 18774 9198 18802 9226
rect 20006 9422 20034 9450
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 13342 8582 13370 8610
rect 13118 8414 13146 8442
rect 13286 8358 13314 8386
rect 20006 8750 20034 8778
rect 18942 8414 18970 8442
rect 20006 8414 20034 8442
rect 18830 8358 18858 8386
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 20006 8105 20034 8106
rect 20006 8079 20007 8105
rect 20007 8079 20033 8105
rect 20033 8079 20034 8105
rect 20006 8078 20034 8079
rect 12670 8022 12698 8050
rect 12166 7742 12194 7770
rect 12782 7769 12810 7770
rect 12782 7743 12783 7769
rect 12783 7743 12809 7769
rect 12809 7743 12810 7769
rect 12782 7742 12810 7743
rect 12950 7713 12978 7714
rect 12950 7687 12951 7713
rect 12951 7687 12977 7713
rect 12977 7687 12978 7713
rect 12950 7686 12978 7687
rect 18830 7686 18858 7714
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 11214 1833 11242 1834
rect 11214 1807 11215 1833
rect 11215 1807 11241 1833
rect 11241 1807 11242 1833
rect 11214 1806 11242 1807
rect 12446 1806 12474 1834
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 13062 1833 13090 1834
rect 13062 1807 13063 1833
rect 13063 1807 13089 1833
rect 13089 1807 13090 1833
rect 13062 1806 13090 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 10761 19110 10766 19138
rect 10794 19110 11214 19138
rect 11242 19110 11247 19138
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 10425 18718 10430 18746
rect 10458 18718 11046 18746
rect 11074 18718 11079 18746
rect 12105 18718 12110 18746
rect 12138 18718 13118 18746
rect 13146 18718 13151 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 11377 13230 11382 13258
rect 11410 13230 11774 13258
rect 11802 13230 12278 13258
rect 12306 13230 12311 13258
rect 9081 13006 9086 13034
rect 9114 13006 9534 13034
rect 9562 13006 9567 13034
rect 9809 13006 9814 13034
rect 9842 13006 10262 13034
rect 10290 13006 10295 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 0 12810 400 12824
rect 0 12782 2086 12810
rect 2114 12782 2119 12810
rect 0 12768 400 12782
rect 10313 12670 10318 12698
rect 10346 12670 10542 12698
rect 10570 12670 11438 12698
rect 11466 12670 13230 12698
rect 13258 12670 13263 12698
rect 7233 12614 7238 12642
rect 7266 12614 8078 12642
rect 8106 12614 8111 12642
rect 8185 12614 8190 12642
rect 8218 12614 10822 12642
rect 10850 12614 12166 12642
rect 12194 12614 12199 12642
rect 12497 12614 12502 12642
rect 12530 12614 13062 12642
rect 13090 12614 13095 12642
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 9585 12446 9590 12474
rect 9618 12446 11046 12474
rect 11074 12446 12054 12474
rect 12082 12446 12087 12474
rect 6897 12390 6902 12418
rect 6930 12390 7630 12418
rect 7658 12390 8134 12418
rect 8162 12390 8862 12418
rect 8890 12390 8895 12418
rect 8353 12334 8358 12362
rect 8386 12334 8806 12362
rect 8834 12334 8839 12362
rect 10369 12334 10374 12362
rect 10402 12334 10934 12362
rect 10962 12334 12614 12362
rect 12642 12334 12647 12362
rect 15946 12334 18830 12362
rect 18858 12334 18863 12362
rect 15946 12306 15974 12334
rect 12217 12278 12222 12306
rect 12250 12278 13006 12306
rect 13034 12278 13039 12306
rect 13169 12278 13174 12306
rect 13202 12278 14070 12306
rect 14098 12278 15974 12306
rect 8913 12222 8918 12250
rect 8946 12222 9590 12250
rect 9618 12222 9814 12250
rect 9842 12222 9847 12250
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 13281 11998 13286 12026
rect 13314 11998 14070 12026
rect 14098 11998 15974 12026
rect 15946 11970 15974 11998
rect 9809 11942 9814 11970
rect 9842 11942 11102 11970
rect 11130 11942 11135 11970
rect 15946 11942 18830 11970
rect 18858 11942 18863 11970
rect 20600 11802 21000 11816
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 8297 11718 8302 11746
rect 8330 11718 8694 11746
rect 8722 11718 8727 11746
rect 12273 11662 12278 11690
rect 12306 11662 12670 11690
rect 12698 11662 12703 11690
rect 8241 11438 8246 11466
rect 8274 11438 8750 11466
rect 8778 11438 8783 11466
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9081 11326 9086 11354
rect 9114 11326 11382 11354
rect 11410 11326 12782 11354
rect 12810 11326 12815 11354
rect 6169 11158 6174 11186
rect 6202 11158 7462 11186
rect 7490 11158 7686 11186
rect 7714 11158 7719 11186
rect 7401 11102 7406 11130
rect 7434 11102 8134 11130
rect 8162 11102 8974 11130
rect 9002 11102 9007 11130
rect 8801 11046 8806 11074
rect 8834 11046 9478 11074
rect 9506 11046 9814 11074
rect 9842 11046 9847 11074
rect 9921 11046 9926 11074
rect 9954 11046 10122 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 7457 10934 7462 10962
rect 7490 10934 9086 10962
rect 9114 10934 9119 10962
rect 10094 10906 10122 11046
rect 8017 10878 8022 10906
rect 8050 10878 8302 10906
rect 8330 10878 8694 10906
rect 8722 10878 8727 10906
rect 9305 10878 9310 10906
rect 9338 10878 10822 10906
rect 10850 10878 10855 10906
rect 11153 10878 11158 10906
rect 11186 10878 13510 10906
rect 13538 10878 14126 10906
rect 14154 10878 14159 10906
rect 10985 10822 10990 10850
rect 11018 10822 12166 10850
rect 12194 10822 12199 10850
rect 2137 10766 2142 10794
rect 2170 10766 6062 10794
rect 6090 10766 6095 10794
rect 12329 10710 12334 10738
rect 12362 10710 15974 10738
rect 15946 10682 15974 10710
rect 15946 10654 18830 10682
rect 18858 10654 18863 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 10929 10486 10934 10514
rect 10962 10486 12614 10514
rect 12642 10486 12726 10514
rect 12754 10486 12759 10514
rect 13393 10486 13398 10514
rect 13426 10486 14182 10514
rect 14210 10486 14215 10514
rect 0 10458 400 10472
rect 20600 10458 21000 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 19945 10430 19950 10458
rect 19978 10430 21000 10458
rect 0 10416 400 10430
rect 20600 10416 21000 10430
rect 6057 10374 6062 10402
rect 6090 10374 6902 10402
rect 6930 10374 6935 10402
rect 10033 10374 10038 10402
rect 10066 10374 11326 10402
rect 11354 10374 11359 10402
rect 7233 10318 7238 10346
rect 7266 10318 7910 10346
rect 7938 10318 10598 10346
rect 10626 10318 10631 10346
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 20600 10122 21000 10136
rect 13449 10094 13454 10122
rect 13482 10094 14182 10122
rect 14210 10094 18942 10122
rect 18970 10094 18975 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 20600 10080 21000 10094
rect 7546 9982 9030 10010
rect 9058 9982 9646 10010
rect 9674 9982 9679 10010
rect 7546 9954 7574 9982
rect 2081 9926 2086 9954
rect 2114 9926 7574 9954
rect 7625 9926 7630 9954
rect 7658 9926 8358 9954
rect 8386 9926 9254 9954
rect 9282 9926 9534 9954
rect 9562 9926 9567 9954
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 7849 9646 7854 9674
rect 7882 9646 8190 9674
rect 8218 9646 8223 9674
rect 8353 9646 8358 9674
rect 8386 9646 9758 9674
rect 9786 9646 9791 9674
rect 10033 9646 10038 9674
rect 10066 9646 12054 9674
rect 12082 9646 12446 9674
rect 12474 9646 13006 9674
rect 13034 9646 13039 9674
rect 2137 9590 2142 9618
rect 2170 9590 6230 9618
rect 6258 9590 8302 9618
rect 8330 9590 8335 9618
rect 9305 9590 9310 9618
rect 9338 9590 9590 9618
rect 9618 9590 9623 9618
rect 11769 9590 11774 9618
rect 11802 9590 12110 9618
rect 12138 9590 12143 9618
rect 8073 9534 8078 9562
rect 8106 9534 9142 9562
rect 9170 9534 9175 9562
rect 9417 9534 9422 9562
rect 9450 9534 10822 9562
rect 10850 9534 11382 9562
rect 11410 9534 11415 9562
rect 7289 9478 7294 9506
rect 7322 9478 7854 9506
rect 7882 9478 7887 9506
rect 9249 9478 9254 9506
rect 9282 9478 9590 9506
rect 9618 9478 9623 9506
rect 10201 9478 10206 9506
rect 10234 9478 10239 9506
rect 10369 9478 10374 9506
rect 10402 9478 10710 9506
rect 10738 9478 11046 9506
rect 11074 9478 11079 9506
rect 11153 9478 11158 9506
rect 11186 9478 12166 9506
rect 12194 9478 12726 9506
rect 12754 9478 12759 9506
rect 14737 9478 14742 9506
rect 14770 9478 18942 9506
rect 18970 9478 18975 9506
rect 0 9450 400 9464
rect 0 9422 966 9450
rect 994 9422 999 9450
rect 0 9408 400 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 8745 9310 8750 9338
rect 8778 9310 9478 9338
rect 9506 9310 9511 9338
rect 9585 9310 9590 9338
rect 9618 9310 10094 9338
rect 10122 9310 10127 9338
rect 10206 9282 10234 9478
rect 20600 9450 21000 9464
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 20600 9408 21000 9422
rect 10761 9310 10766 9338
rect 10794 9310 11886 9338
rect 11914 9310 11919 9338
rect 15946 9310 18830 9338
rect 18858 9310 18863 9338
rect 15946 9282 15974 9310
rect 7401 9254 7406 9282
rect 7434 9254 9030 9282
rect 9058 9254 9646 9282
rect 9674 9254 9926 9282
rect 9954 9254 10234 9282
rect 10593 9254 10598 9282
rect 10626 9254 10822 9282
rect 10850 9254 11214 9282
rect 11242 9254 11247 9282
rect 14345 9254 14350 9282
rect 14378 9254 14630 9282
rect 14658 9254 15974 9282
rect 7009 9198 7014 9226
rect 7042 9198 7686 9226
rect 7714 9198 9254 9226
rect 9282 9198 9287 9226
rect 9473 9198 9478 9226
rect 9506 9198 9702 9226
rect 9730 9198 10094 9226
rect 10122 9198 10127 9226
rect 14457 9198 14462 9226
rect 14490 9198 18774 9226
rect 18802 9198 18807 9226
rect 7961 9142 7966 9170
rect 7994 9142 8862 9170
rect 8890 9142 8895 9170
rect 20600 9114 21000 9128
rect 9865 9086 9870 9114
rect 9898 9086 10206 9114
rect 10234 9086 10239 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 8801 8862 8806 8890
rect 8834 8862 9086 8890
rect 9114 8862 9119 8890
rect 8409 8806 8414 8834
rect 8442 8806 8918 8834
rect 8946 8806 9198 8834
rect 9226 8806 9310 8834
rect 9338 8806 9343 8834
rect 9473 8806 9478 8834
rect 9506 8806 9926 8834
rect 9954 8806 10878 8834
rect 10906 8806 12054 8834
rect 12082 8806 12087 8834
rect 12329 8806 12334 8834
rect 12362 8806 12614 8834
rect 12642 8806 12647 8834
rect 20600 8778 21000 8792
rect 9753 8750 9758 8778
rect 9786 8750 10654 8778
rect 10682 8750 10687 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 7345 8694 7350 8722
rect 7378 8694 9702 8722
rect 9730 8694 9735 8722
rect 11769 8694 11774 8722
rect 11802 8694 12110 8722
rect 12138 8694 12143 8722
rect 12721 8694 12726 8722
rect 12754 8694 13118 8722
rect 13146 8694 13151 8722
rect 8913 8638 8918 8666
rect 8946 8638 9590 8666
rect 9618 8638 9623 8666
rect 10089 8638 10094 8666
rect 10122 8638 10141 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 2137 8582 2142 8610
rect 2170 8582 7294 8610
rect 7322 8582 8358 8610
rect 8386 8582 8391 8610
rect 10257 8582 10262 8610
rect 10290 8582 10654 8610
rect 10682 8582 11102 8610
rect 11130 8582 11135 8610
rect 11601 8582 11606 8610
rect 11634 8582 13342 8610
rect 13370 8582 13375 8610
rect 11606 8554 11634 8582
rect 9977 8526 9982 8554
rect 10010 8526 10318 8554
rect 10346 8526 11634 8554
rect 7121 8470 7126 8498
rect 7154 8470 8750 8498
rect 8778 8470 8783 8498
rect 10929 8470 10934 8498
rect 10962 8470 11494 8498
rect 11522 8470 11886 8498
rect 11914 8470 11919 8498
rect 12217 8470 12222 8498
rect 12250 8470 12558 8498
rect 12586 8470 12591 8498
rect 20600 8442 21000 8456
rect 8353 8414 8358 8442
rect 8386 8414 8638 8442
rect 8666 8414 8671 8442
rect 9697 8414 9702 8442
rect 9730 8414 9926 8442
rect 9954 8414 10150 8442
rect 10178 8414 10183 8442
rect 10761 8414 10766 8442
rect 10794 8414 11998 8442
rect 12026 8414 12031 8442
rect 13113 8414 13118 8442
rect 13146 8414 18942 8442
rect 18970 8414 18975 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 20600 8400 21000 8414
rect 11657 8358 11662 8386
rect 11690 8358 12054 8386
rect 12082 8358 12087 8386
rect 13281 8358 13286 8386
rect 13314 8358 18830 8386
rect 18858 8358 18863 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 0 8106 400 8120
rect 20600 8106 21000 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 20001 8078 20006 8106
rect 20034 8078 21000 8106
rect 0 8064 400 8078
rect 20600 8064 21000 8078
rect 8465 8022 8470 8050
rect 8498 8022 9814 8050
rect 9842 8022 10094 8050
rect 10122 8022 10127 8050
rect 11769 8022 11774 8050
rect 11802 8022 12670 8050
rect 12698 8022 12703 8050
rect 10089 7966 10094 7994
rect 10122 7966 10598 7994
rect 10626 7966 10631 7994
rect 9529 7910 9534 7938
rect 9562 7910 10038 7938
rect 10066 7910 10990 7938
rect 11018 7910 11023 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 12161 7742 12166 7770
rect 12194 7742 12782 7770
rect 12810 7742 12815 7770
rect 7457 7686 7462 7714
rect 7490 7686 7854 7714
rect 7882 7686 7887 7714
rect 12945 7686 12950 7714
rect 12978 7686 18830 7714
rect 18858 7686 18863 7714
rect 7289 7630 7294 7658
rect 7322 7630 7798 7658
rect 7826 7630 8414 7658
rect 8442 7630 8447 7658
rect 10929 7574 10934 7602
rect 10962 7574 11718 7602
rect 11746 7574 11751 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 9529 6678 9534 6706
rect 9562 6678 10206 6706
rect 10234 6678 10239 6706
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 7737 2590 7742 2618
rect 7770 2590 8358 2618
rect 8386 2590 8391 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 10089 2030 10094 2058
rect 10122 2030 10710 2058
rect 10738 2030 10743 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10761 1806 10766 1834
rect 10794 1806 11214 1834
rect 11242 1806 11247 1834
rect 12441 1806 12446 1834
rect 12474 1806 13062 1834
rect 13090 1806 13095 1834
rect 8073 1694 8078 1722
rect 8106 1694 9254 1722
rect 9282 1694 9287 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 10094 8638 10122 8666
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 10094 8022 10122 8050
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 10094 8666 10122 8671
rect 10094 8050 10122 8638
rect 10094 8017 10122 8022
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _068_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11536 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _069_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10752 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _070_
timestamp 1698175906
transform -1 0 10416 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _071_
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _072_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12432 0 1 8624
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _073_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12264 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _074_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _075_
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _076_
timestamp 1698175906
transform 1 0 11984 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _077_
timestamp 1698175906
transform -1 0 11816 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _078_
timestamp 1698175906
transform -1 0 13608 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _079_
timestamp 1698175906
transform -1 0 13216 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _080_
timestamp 1698175906
transform -1 0 10864 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _081_
timestamp 1698175906
transform 1 0 9744 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _082_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7616 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _083_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _084_
timestamp 1698175906
transform 1 0 8848 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _085_
timestamp 1698175906
transform -1 0 11200 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _086_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _087_
timestamp 1698175906
transform -1 0 9016 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _088_
timestamp 1698175906
transform -1 0 9800 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _089_
timestamp 1698175906
transform -1 0 10192 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _090_
timestamp 1698175906
transform 1 0 9240 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _091_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10920 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _092_
timestamp 1698175906
transform 1 0 10920 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _093_
timestamp 1698175906
transform -1 0 12152 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _094_
timestamp 1698175906
transform 1 0 11200 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _095_
timestamp 1698175906
transform 1 0 10920 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10248 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _097_
timestamp 1698175906
transform -1 0 9576 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7616 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _099_
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10136 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _101_
timestamp 1698175906
transform 1 0 11984 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _102_
timestamp 1698175906
transform -1 0 11480 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_
timestamp 1698175906
transform -1 0 10920 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7952 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10752 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9016 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10976 0 -1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _109_
timestamp 1698175906
transform 1 0 11536 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1698175906
transform 1 0 8176 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _111_
timestamp 1698175906
transform -1 0 8344 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform 1 0 8680 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_
timestamp 1698175906
transform 1 0 10024 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _114_
timestamp 1698175906
transform 1 0 10080 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _115_
timestamp 1698175906
transform 1 0 9632 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _116_
timestamp 1698175906
transform 1 0 9576 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _117_
timestamp 1698175906
transform 1 0 7784 0 -1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _118_
timestamp 1698175906
transform 1 0 6832 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7056 0 1 10192
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _120_
timestamp 1698175906
transform -1 0 9688 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _121_
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_
timestamp 1698175906
transform 1 0 14056 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_
timestamp 1698175906
transform -1 0 13496 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 12880 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 10808 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1698175906
transform -1 0 13328 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _127_
timestamp 1698175906
transform 1 0 12096 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _128_
timestamp 1698175906
transform -1 0 8344 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 8456 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform -1 0 9408 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _131_
timestamp 1698175906
transform 1 0 7728 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform 1 0 13160 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _133_
timestamp 1698175906
transform 1 0 12600 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform -1 0 8568 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _135_
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _137_
timestamp 1698175906
transform 1 0 10808 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _138_
timestamp 1698175906
transform -1 0 7728 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _139_
timestamp 1698175906
transform 1 0 6776 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _140_
timestamp 1698175906
transform 1 0 9128 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _141_
timestamp 1698175906
transform 1 0 6888 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _142_
timestamp 1698175906
transform -1 0 7616 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _143_
timestamp 1698175906
transform 1 0 8008 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _145_
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _146_
timestamp 1698175906
transform -1 0 7784 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _147_
timestamp 1698175906
transform 1 0 12544 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _148_
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _149_
timestamp 1698175906
transform 1 0 10248 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _150_
timestamp 1698175906
transform 1 0 8792 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _151_
timestamp 1698175906
transform 1 0 11648 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _152_
timestamp 1698175906
transform -1 0 11088 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _153_
timestamp 1698175906
transform 1 0 11592 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _154_
timestamp 1698175906
transform 1 0 12656 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _155_
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform -1 0 7896 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 7224 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _161_
timestamp 1698175906
transform 1 0 13048 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform -1 0 11088 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _163_
timestamp 1698175906
transform 1 0 12712 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _164_
timestamp 1698175906
transform 1 0 14224 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform 1 0 7896 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9016 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9576 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11256 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout25
timestamp 1698175906
transform 1 0 8008 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_52 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3584 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_60 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4032 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_65 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698175906
transform 1 0 4424 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_104 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_108
timestamp 1698175906
transform 1 0 6720 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_164
timestamp 1698175906
transform 1 0 9856 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_168
timestamp 1698175906
transform 1 0 10080 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_210
timestamp 1698175906
transform 1 0 12432 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 13944 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_256
timestamp 1698175906
transform 1 0 15008 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_258
timestamp 1698175906
transform 1 0 15120 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_263
timestamp 1698175906
transform 1 0 15400 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698175906
transform 1 0 15848 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_158
timestamp 1698175906
transform 1 0 9520 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_166
timestamp 1698175906
transform 1 0 9968 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_168
timestamp 1698175906
transform 1 0 10080 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195
timestamp 1698175906
transform 1 0 11592 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 12040 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_123
timestamp 1698175906
transform 1 0 7560 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_153
timestamp 1698175906
transform 1 0 9240 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_169
timestamp 1698175906
transform 1 0 10136 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_173
timestamp 1698175906
transform 1 0 10360 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698175906
transform 1 0 9072 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_154
timestamp 1698175906
transform 1 0 9296 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_156
timestamp 1698175906
transform 1 0 9408 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_186
timestamp 1698175906
transform 1 0 11088 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_202
timestamp 1698175906
transform 1 0 11984 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_193
timestamp 1698175906
transform 1 0 11480 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_224
timestamp 1698175906
transform 1 0 13216 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 14112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_112
timestamp 1698175906
transform 1 0 6944 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_116
timestamp 1698175906
transform 1 0 7168 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_135
timestamp 1698175906
transform 1 0 8232 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 8456 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_150
timestamp 1698175906
transform 1 0 9072 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_186
timestamp 1698175906
transform 1 0 11088 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_202
timestamp 1698175906
transform 1 0 11984 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_221
timestamp 1698175906
transform 1 0 13048 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_253
timestamp 1698175906
transform 1 0 14840 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_269
timestamp 1698175906
transform 1 0 15736 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_141
timestamp 1698175906
transform 1 0 8568 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_157
timestamp 1698175906
transform 1 0 9464 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_161
timestamp 1698175906
transform 1 0 9688 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_185
timestamp 1698175906
transform 1 0 11032 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_193
timestamp 1698175906
transform 1 0 11480 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_195
timestamp 1698175906
transform 1 0 11592 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_225
timestamp 1698175906
transform 1 0 13272 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698175906
transform 1 0 6720 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698175906
transform 1 0 6832 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_150
timestamp 1698175906
transform 1 0 9072 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_158
timestamp 1698175906
transform 1 0 9520 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_173
timestamp 1698175906
transform 1 0 10360 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_189
timestamp 1698175906
transform 1 0 11256 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_220
timestamp 1698175906
transform 1 0 12992 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_227
timestamp 1698175906
transform 1 0 13384 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_259
timestamp 1698175906
transform 1 0 15176 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 16072 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_139
timestamp 1698175906
transform 1 0 8456 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 10360 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_183
timestamp 1698175906
transform 1 0 10920 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_199
timestamp 1698175906
transform 1 0 11816 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_201
timestamp 1698175906
transform 1 0 11928 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_217
timestamp 1698175906
transform 1 0 12824 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_233
timestamp 1698175906
transform 1 0 13720 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 14168 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_96
timestamp 1698175906
transform 1 0 6048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_127
timestamp 1698175906
transform 1 0 7784 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 8232 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_149
timestamp 1698175906
transform 1 0 9016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_157
timestamp 1698175906
transform 1 0 9464 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_188
timestamp 1698175906
transform 1 0 11200 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_204
timestamp 1698175906
transform 1 0 12096 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_218
timestamp 1698175906
transform 1 0 12880 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_222
timestamp 1698175906
transform 1 0 13104 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_229
timestamp 1698175906
transform 1 0 13496 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_237
timestamp 1698175906
transform 1 0 13944 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_241
timestamp 1698175906
transform 1 0 14168 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_248
timestamp 1698175906
transform 1 0 14560 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_125
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_139
timestamp 1698175906
transform 1 0 8456 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_147
timestamp 1698175906
transform 1 0 8904 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_193
timestamp 1698175906
transform 1 0 11480 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_209
timestamp 1698175906
transform 1 0 12376 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_213
timestamp 1698175906
transform 1 0 12600 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_253
timestamp 1698175906
transform 1 0 14840 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_285
timestamp 1698175906
transform 1 0 16632 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_301
timestamp 1698175906
transform 1 0 17528 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_309
timestamp 1698175906
transform 1 0 17976 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_313
timestamp 1698175906
transform 1 0 18200 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_92
timestamp 1698175906
transform 1 0 5824 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_94
timestamp 1698175906
transform 1 0 5936 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_124
timestamp 1698175906
transform 1 0 7616 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_126
timestamp 1698175906
transform 1 0 7728 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698175906
transform 1 0 8848 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_148
timestamp 1698175906
transform 1 0 8960 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_243
timestamp 1698175906
transform 1 0 14280 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698175906
transform 1 0 16072 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 16296 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698175906
transform 1 0 6776 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698175906
transform 1 0 10696 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_188
timestamp 1698175906
transform 1 0 11200 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_96
timestamp 1698175906
transform 1 0 6048 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_126
timestamp 1698175906
transform 1 0 7728 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698175906
transform 1 0 8344 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 8456 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698175906
transform 1 0 9072 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698175906
transform 1 0 12768 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_218
timestamp 1698175906
transform 1 0 12880 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_224
timestamp 1698175906
transform 1 0 13216 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_231
timestamp 1698175906
transform 1 0 13608 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_263
timestamp 1698175906
transform 1 0 15400 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 7112 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_117
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_139
timestamp 1698175906
transform 1 0 8456 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_151
timestamp 1698175906
transform 1 0 9128 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_159
timestamp 1698175906
transform 1 0 9576 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_161
timestamp 1698175906
transform 1 0 9688 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_170
timestamp 1698175906
transform 1 0 10192 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_182
timestamp 1698175906
transform 1 0 10864 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_189
timestamp 1698175906
transform 1 0 11256 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_221
timestamp 1698175906
transform 1 0 13048 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_237
timestamp 1698175906
transform 1 0 13944 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_104
timestamp 1698175906
transform 1 0 6496 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_120
timestamp 1698175906
transform 1 0 7392 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_128
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_132
timestamp 1698175906
transform 1 0 8064 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_146
timestamp 1698175906
transform 1 0 8848 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_162
timestamp 1698175906
transform 1 0 9744 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_170
timestamp 1698175906
transform 1 0 10192 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_174
timestamp 1698175906
transform 1 0 10416 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_181
timestamp 1698175906
transform 1 0 10808 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_197
timestamp 1698175906
transform 1 0 11704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 12152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_221
timestamp 1698175906
transform 1 0 13048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_228
timestamp 1698175906
transform 1 0 13440 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_260
timestamp 1698175906
transform 1 0 15232 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698175906
transform 1 0 7560 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_160
timestamp 1698175906
transform 1 0 9632 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698175906
transform 1 0 10080 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 10304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698175906
transform 1 0 11032 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698175906
transform 1 0 11144 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_196
timestamp 1698175906
transform 1 0 11648 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_104
timestamp 1698175906
transform 1 0 6496 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_108
timestamp 1698175906
transform 1 0 6720 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_152
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_164
timestamp 1698175906
transform 1 0 9856 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_168
timestamp 1698175906
transform 1 0 10080 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_170
timestamp 1698175906
transform 1 0 10192 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698175906
transform 1 0 12152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_241
timestamp 1698175906
transform 1 0 14168 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 15960 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 16184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_131
timestamp 1698175906
transform 1 0 8008 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_137
timestamp 1698175906
transform 1 0 8344 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_210
timestamp 1698175906
transform 1 0 12432 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_218
timestamp 1698175906
transform 1 0 12880 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_220
timestamp 1698175906
transform 1 0 12992 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_226
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_150
timestamp 1698175906
transform 1 0 9072 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_154
timestamp 1698175906
transform 1 0 9296 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_161
timestamp 1698175906
transform 1 0 9688 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_174
timestamp 1698175906
transform 1 0 10416 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_178
timestamp 1698175906
transform 1 0 10640 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_188
timestamp 1698175906
transform 1 0 11200 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_194
timestamp 1698175906
transform 1 0 11536 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 16128 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 14168 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_174
timestamp 1698175906
transform 1 0 10416 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 11928 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita14_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4312 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita14_27
timestamp 1698175906
transform -1 0 15400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 12488 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 8288 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 7784 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 10136 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 10472 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 4032 0 4088 400 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 7392 0 7448 400 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 15120 0 15176 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 7728 0 7784 400 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 9408 400 9464 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 8064 0 8120 400 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 11312 12012 11312 12012 0 _000_
rlabel metal2 11676 10192 11676 10192 0 _001_
rlabel metal2 7420 11172 7420 11172 0 _002_
rlabel metal2 7252 12516 7252 12516 0 _003_
rlabel metal2 9688 7700 9688 7700 0 _004_
rlabel metal2 7364 8596 7364 8596 0 _005_
rlabel metal2 7252 10164 7252 10164 0 _006_
rlabel metal2 8484 12068 8484 12068 0 _007_
rlabel metal2 13244 9436 13244 9436 0 _008_
rlabel metal2 12236 12152 12236 12152 0 _009_
rlabel metal2 7308 9352 7308 9352 0 _010_
rlabel metal2 12740 11788 12740 11788 0 _011_
rlabel metal2 7140 8288 7140 8288 0 _012_
rlabel metal2 10808 12404 10808 12404 0 _013_
rlabel metal2 9548 12572 9548 12572 0 _014_
rlabel metal2 12124 8232 12124 8232 0 _015_
rlabel metal2 10668 6916 10668 6916 0 _016_
rlabel metal3 11872 8372 11872 8372 0 _017_
rlabel metal2 13104 10052 13104 10052 0 _018_
rlabel metal2 9660 11004 9660 11004 0 _019_
rlabel metal2 10612 8008 10612 8008 0 _020_
rlabel metal2 11788 8568 11788 8568 0 _021_
rlabel metal2 13244 10780 13244 10780 0 _022_
rlabel metal2 10388 11172 10388 11172 0 _023_
rlabel metal2 8260 11228 8260 11228 0 _024_
rlabel metal2 7476 10696 7476 10696 0 _025_
rlabel metal3 10556 9492 10556 9492 0 _026_
rlabel metal3 8540 9268 8540 9268 0 _027_
rlabel metal3 9156 8036 9156 8036 0 _028_
rlabel metal2 10332 9324 10332 9324 0 _029_
rlabel metal2 11284 11928 11284 11928 0 _030_
rlabel metal2 9408 9268 9408 9268 0 _031_
rlabel metal2 10780 10388 10780 10388 0 _032_
rlabel metal2 13524 10864 13524 10864 0 _033_
rlabel metal2 11620 11984 11620 11984 0 _034_
rlabel metal3 11676 9492 11676 9492 0 _035_
rlabel via2 8372 9660 8372 9660 0 _036_
rlabel metal3 9408 9940 9408 9940 0 _037_
rlabel metal2 8708 10920 8708 10920 0 _038_
rlabel metal2 9828 10584 9828 10584 0 _039_
rlabel metal2 12068 9632 12068 9632 0 _040_
rlabel metal3 11956 9604 11956 9604 0 _041_
rlabel metal2 10612 9240 10612 9240 0 _042_
rlabel metal2 10836 10668 10836 10668 0 _043_
rlabel metal2 8148 11508 8148 11508 0 _044_
rlabel metal2 11564 9744 11564 9744 0 _045_
rlabel metal2 9100 9744 9100 9744 0 _046_
rlabel metal2 10892 9016 10892 9016 0 _047_
rlabel metal2 11900 9016 11900 9016 0 _048_
rlabel metal2 8316 12684 8316 12684 0 _049_
rlabel metal2 9604 8736 9604 8736 0 _050_
rlabel metal2 10192 8540 10192 8540 0 _051_
rlabel metal2 11620 8512 11620 8512 0 _052_
rlabel metal2 7924 10220 7924 10220 0 _053_
rlabel metal2 7028 10388 7028 10388 0 _054_
rlabel metal2 9100 12684 9100 12684 0 _055_
rlabel metal2 13412 9884 13412 9884 0 _056_
rlabel metal3 12488 11676 12488 11676 0 _057_
rlabel metal2 13244 12152 13244 12152 0 _058_
rlabel metal2 12516 12292 12516 12292 0 _059_
rlabel metal2 7980 9352 7980 9352 0 _060_
rlabel metal2 7812 9632 7812 9632 0 _061_
rlabel metal3 8624 9548 8624 9548 0 _062_
rlabel metal2 13020 11508 13020 11508 0 _063_
rlabel metal2 8344 8036 8344 8036 0 _064_
rlabel metal2 11228 13132 11228 13132 0 _065_
rlabel metal2 9828 12684 9828 12684 0 _066_
rlabel metal2 12236 8456 12236 8456 0 _067_
rlabel metal3 1239 12796 1239 12796 0 clk
rlabel metal2 11340 10220 11340 10220 0 clknet_0_clk
rlabel metal2 6916 12376 6916 12376 0 clknet_1_0__leaf_clk
rlabel metal3 11340 7588 11340 7588 0 clknet_1_1__leaf_clk
rlabel metal3 6832 11172 6832 11172 0 dut14.count\[0\]
rlabel metal2 8708 11676 8708 11676 0 dut14.count\[1\]
rlabel metal2 11116 8876 11116 8876 0 dut14.count\[2\]
rlabel metal3 8820 8820 8820 8820 0 dut14.count\[3\]
rlabel metal2 8176 8092 8176 8092 0 net1
rlabel metal2 18956 8624 18956 8624 0 net10
rlabel metal2 10836 4732 10836 4732 0 net11
rlabel metal2 10220 4424 10220 4424 0 net12
rlabel metal3 15022 12012 15022 12012 0 net13
rlabel metal3 11844 13244 11844 13244 0 net14
rlabel metal2 10416 15960 10416 15960 0 net15
rlabel metal2 6244 9380 6244 9380 0 net16
rlabel metal3 15022 12292 15022 12292 0 net17
rlabel metal2 14476 9240 14476 9240 0 net18
rlabel metal3 6496 10388 6496 10388 0 net19
rlabel metal2 18844 7868 18844 7868 0 net2
rlabel metal2 8316 1764 8316 1764 0 net20
rlabel metal3 15960 10696 15960 10696 0 net21
rlabel metal2 10696 15960 10696 15960 0 net22
rlabel metal2 12628 16030 12628 16030 0 net23
rlabel metal2 9716 19012 9716 19012 0 net24
rlabel metal2 2156 8512 2156 8512 0 net25
rlabel metal2 4060 1015 4060 1015 0 net26
rlabel metal2 15148 1015 15148 1015 0 net27
rlabel metal2 12628 2982 12628 2982 0 net3
rlabel metal2 13468 10472 13468 10472 0 net4
rlabel metal2 7812 7812 7812 7812 0 net5
rlabel metal2 18956 9352 18956 9352 0 net6
rlabel metal3 7672 7700 7672 7700 0 net7
rlabel metal2 14224 10276 14224 10276 0 net8
rlabel metal2 18844 8400 18844 8400 0 net9
rlabel metal3 679 8092 679 8092 0 segm[10]
rlabel metal3 20321 8092 20321 8092 0 segm[11]
rlabel metal2 12460 1099 12460 1099 0 segm[12]
rlabel metal2 19964 10584 19964 10584 0 segm[13]
rlabel metal2 7420 1043 7420 1043 0 segm[1]
rlabel metal3 20321 9100 20321 9100 0 segm[2]
rlabel metal2 7756 1491 7756 1491 0 segm[4]
rlabel metal2 20020 9548 20020 9548 0 segm[5]
rlabel metal2 20020 8400 20020 8400 0 segm[6]
rlabel metal2 20020 8820 20020 8820 0 segm[7]
rlabel metal2 10780 1099 10780 1099 0 segm[8]
rlabel metal2 10108 1211 10108 1211 0 segm[9]
rlabel metal2 20020 11900 20020 11900 0 sel[0]
rlabel metal2 11788 19873 11788 19873 0 sel[10]
rlabel metal2 10444 19677 10444 19677 0 sel[11]
rlabel metal3 679 9436 679 9436 0 sel[1]
rlabel metal2 20020 12180 20020 12180 0 sel[2]
rlabel metal2 20020 9828 20020 9828 0 sel[3]
rlabel metal3 679 10444 679 10444 0 sel[4]
rlabel metal2 8092 1043 8092 1043 0 sel[5]
rlabel metal2 20020 10276 20020 10276 0 sel[6]
rlabel metal2 10780 19873 10780 19873 0 sel[7]
rlabel metal2 12124 19677 12124 19677 0 sel[8]
rlabel metal2 9436 19845 9436 19845 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
