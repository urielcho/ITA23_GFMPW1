magic
tech gf180mcuD
magscale 1 5
timestamp 1699642983
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 14687 19137 14713 19143
rect 14687 19105 14713 19111
rect 9025 18999 9031 19025
rect 9057 18999 9063 19025
rect 10705 18999 10711 19025
rect 10737 18999 10743 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 14289 18999 14295 19025
rect 14321 18999 14327 19025
rect 8639 18969 8665 18975
rect 8639 18937 8665 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 13119 18745 13145 18751
rect 13119 18713 13145 18719
rect 14575 18745 14601 18751
rect 14575 18713 14601 18719
rect 12609 18607 12615 18633
rect 12641 18607 12647 18633
rect 14065 18607 14071 18633
rect 14097 18607 14103 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 855 18185 881 18191
rect 855 18153 881 18159
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 12217 14351 12223 14377
rect 12249 14351 12255 14377
rect 12391 14321 12417 14327
rect 10817 14295 10823 14321
rect 10849 14295 10855 14321
rect 12391 14289 12417 14295
rect 12783 14265 12809 14271
rect 11153 14239 11159 14265
rect 11185 14239 11191 14265
rect 12553 14239 12559 14265
rect 12585 14239 12591 14265
rect 12783 14233 12809 14239
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 11159 14041 11185 14047
rect 11159 14009 11185 14015
rect 12279 14041 12305 14047
rect 12279 14009 12305 14015
rect 11103 13929 11129 13935
rect 2137 13903 2143 13929
rect 2169 13903 2175 13929
rect 9305 13903 9311 13929
rect 9337 13903 9343 13929
rect 11103 13897 11129 13903
rect 11215 13929 11241 13935
rect 11215 13897 11241 13903
rect 11439 13929 11465 13935
rect 11439 13897 11465 13903
rect 12167 13929 12193 13935
rect 12167 13897 12193 13903
rect 12335 13929 12361 13935
rect 12609 13903 12615 13929
rect 12641 13903 12647 13929
rect 12335 13897 12361 13903
rect 10991 13873 11017 13879
rect 14295 13873 14321 13879
rect 9641 13847 9647 13873
rect 9673 13847 9679 13873
rect 10705 13847 10711 13873
rect 10737 13847 10743 13873
rect 13001 13847 13007 13873
rect 13033 13847 13039 13873
rect 14065 13847 14071 13873
rect 14097 13847 14103 13873
rect 10991 13841 11017 13847
rect 14295 13841 14321 13847
rect 967 13817 993 13823
rect 967 13785 993 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 12111 13593 12137 13599
rect 1017 13567 1023 13593
rect 1049 13567 1055 13593
rect 13785 13567 13791 13593
rect 13817 13567 13823 13593
rect 12111 13561 12137 13567
rect 12055 13537 12081 13543
rect 14015 13537 14041 13543
rect 2137 13511 2143 13537
rect 2169 13511 2175 13537
rect 12385 13511 12391 13537
rect 12417 13511 12423 13537
rect 12055 13505 12081 13511
rect 14015 13505 14041 13511
rect 7463 13481 7489 13487
rect 7289 13455 7295 13481
rect 7321 13455 7327 13481
rect 7463 13449 7489 13455
rect 9983 13481 10009 13487
rect 9983 13449 10009 13455
rect 10151 13481 10177 13487
rect 12721 13455 12727 13481
rect 12753 13455 12759 13481
rect 10151 13449 10177 13455
rect 11943 13425 11969 13431
rect 11943 13393 11969 13399
rect 12167 13425 12193 13431
rect 12167 13393 12193 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8919 13257 8945 13263
rect 7625 13231 7631 13257
rect 7657 13231 7663 13257
rect 8919 13225 8945 13231
rect 9143 13257 9169 13263
rect 9143 13225 9169 13231
rect 9255 13257 9281 13263
rect 9255 13225 9281 13231
rect 10487 13257 10513 13263
rect 10487 13225 10513 13231
rect 12671 13257 12697 13263
rect 12671 13225 12697 13231
rect 12727 13257 12753 13263
rect 12727 13225 12753 13231
rect 13119 13257 13145 13263
rect 13119 13225 13145 13231
rect 13231 13257 13257 13263
rect 13231 13225 13257 13231
rect 13511 13257 13537 13263
rect 13511 13225 13537 13231
rect 13287 13201 13313 13207
rect 13287 13169 13313 13175
rect 13567 13201 13593 13207
rect 13567 13169 13593 13175
rect 8807 13145 8833 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 7401 13119 7407 13145
rect 7433 13119 7439 13145
rect 7737 13119 7743 13145
rect 7769 13119 7775 13145
rect 8689 13119 8695 13145
rect 8721 13119 8727 13145
rect 8807 13113 8833 13119
rect 8975 13145 9001 13151
rect 8975 13113 9001 13119
rect 9311 13145 9337 13151
rect 9311 13113 9337 13119
rect 10431 13145 10457 13151
rect 10431 13113 10457 13119
rect 10599 13145 10625 13151
rect 10599 13113 10625 13119
rect 10711 13145 10737 13151
rect 10711 13113 10737 13119
rect 12615 13145 12641 13151
rect 12615 13113 12641 13119
rect 12951 13145 12977 13151
rect 12951 13113 12977 13119
rect 13399 13145 13425 13151
rect 13399 13113 13425 13119
rect 8023 13089 8049 13095
rect 5945 13063 5951 13089
rect 5977 13063 5983 13089
rect 7065 13063 7071 13089
rect 7097 13063 7103 13089
rect 8745 13063 8751 13089
rect 8777 13063 8783 13089
rect 8023 13057 8049 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 6903 12865 6929 12871
rect 6903 12833 6929 12839
rect 9255 12809 9281 12815
rect 7961 12783 7967 12809
rect 7993 12783 7999 12809
rect 9025 12783 9031 12809
rect 9057 12783 9063 12809
rect 9255 12777 9281 12783
rect 11887 12809 11913 12815
rect 11887 12777 11913 12783
rect 12167 12809 12193 12815
rect 12167 12777 12193 12783
rect 20007 12809 20033 12815
rect 20007 12777 20033 12783
rect 10095 12753 10121 12759
rect 7625 12727 7631 12753
rect 7657 12727 7663 12753
rect 10095 12721 10121 12727
rect 10207 12753 10233 12759
rect 11663 12753 11689 12759
rect 10369 12727 10375 12753
rect 10401 12727 10407 12753
rect 10929 12727 10935 12753
rect 10961 12727 10967 12753
rect 11153 12727 11159 12753
rect 11185 12727 11191 12753
rect 10207 12721 10233 12727
rect 11663 12721 11689 12727
rect 11943 12753 11969 12759
rect 11943 12721 11969 12727
rect 12055 12753 12081 12759
rect 12055 12721 12081 12727
rect 12223 12753 12249 12759
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 12223 12721 12249 12727
rect 6959 12697 6985 12703
rect 11775 12697 11801 12703
rect 10649 12671 10655 12697
rect 10681 12671 10687 12697
rect 11433 12671 11439 12697
rect 11465 12671 11471 12697
rect 6959 12665 6985 12671
rect 11775 12665 11801 12671
rect 12391 12697 12417 12703
rect 12391 12665 12417 12671
rect 10705 12615 10711 12641
rect 10737 12615 10743 12641
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7239 12473 7265 12479
rect 7239 12441 7265 12447
rect 7743 12473 7769 12479
rect 7743 12441 7769 12447
rect 7799 12473 7825 12479
rect 11271 12473 11297 12479
rect 8857 12447 8863 12473
rect 8889 12447 8895 12473
rect 9137 12447 9143 12473
rect 9169 12447 9175 12473
rect 7799 12441 7825 12447
rect 11271 12441 11297 12447
rect 11663 12473 11689 12479
rect 14911 12473 14937 12479
rect 12889 12447 12895 12473
rect 12921 12447 12927 12473
rect 11663 12441 11689 12447
rect 14911 12441 14937 12447
rect 7575 12417 7601 12423
rect 9865 12391 9871 12417
rect 9897 12391 9903 12417
rect 7575 12385 7601 12391
rect 7687 12361 7713 12367
rect 8695 12361 8721 12367
rect 11439 12361 11465 12367
rect 7009 12335 7015 12361
rect 7041 12335 7047 12361
rect 7905 12335 7911 12361
rect 7937 12335 7943 12361
rect 9249 12335 9255 12361
rect 9281 12335 9287 12361
rect 9473 12335 9479 12361
rect 9505 12335 9511 12361
rect 7687 12329 7713 12335
rect 8695 12329 8721 12335
rect 11439 12329 11465 12335
rect 13063 12361 13089 12367
rect 13225 12335 13231 12361
rect 13257 12335 13263 12361
rect 13063 12329 13089 12335
rect 5553 12279 5559 12305
rect 5585 12279 5591 12305
rect 6617 12279 6623 12305
rect 6649 12279 6655 12305
rect 10929 12279 10935 12305
rect 10961 12279 10967 12305
rect 13617 12279 13623 12305
rect 13649 12279 13655 12305
rect 14681 12279 14687 12305
rect 14713 12279 14719 12305
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 13847 12081 13873 12087
rect 13847 12049 13873 12055
rect 967 12025 993 12031
rect 11495 12025 11521 12031
rect 11265 11999 11271 12025
rect 11297 11999 11303 12025
rect 967 11993 993 11999
rect 11495 11993 11521 11999
rect 13399 12025 13425 12031
rect 13399 11993 13425 11999
rect 13679 11969 13705 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 11153 11943 11159 11969
rect 11185 11943 11191 11969
rect 13679 11937 13705 11943
rect 13791 11969 13817 11975
rect 13791 11937 13817 11943
rect 6847 11913 6873 11919
rect 6847 11881 6873 11887
rect 6903 11913 6929 11919
rect 8191 11913 8217 11919
rect 7737 11887 7743 11913
rect 7769 11887 7775 11913
rect 6903 11881 6929 11887
rect 8191 11881 8217 11887
rect 13847 11913 13873 11919
rect 13847 11881 13873 11887
rect 6735 11857 6761 11863
rect 6735 11825 6761 11831
rect 7911 11857 7937 11863
rect 7911 11825 7937 11831
rect 8023 11857 8049 11863
rect 8023 11825 8049 11831
rect 8135 11857 8161 11863
rect 8135 11825 8161 11831
rect 13343 11857 13369 11863
rect 13343 11825 13369 11831
rect 13455 11857 13481 11863
rect 13455 11825 13481 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 6511 11689 6537 11695
rect 6511 11657 6537 11663
rect 6623 11689 6649 11695
rect 6623 11657 6649 11663
rect 8639 11689 8665 11695
rect 8639 11657 8665 11663
rect 8751 11689 8777 11695
rect 14407 11689 14433 11695
rect 9305 11663 9311 11689
rect 9337 11663 9343 11689
rect 8751 11657 8777 11663
rect 14407 11657 14433 11663
rect 6679 11633 6705 11639
rect 12167 11633 12193 11639
rect 7233 11607 7239 11633
rect 7265 11607 7271 11633
rect 11041 11607 11047 11633
rect 11073 11607 11079 11633
rect 11769 11607 11775 11633
rect 11801 11607 11807 11633
rect 6679 11601 6705 11607
rect 12167 11601 12193 11607
rect 8807 11577 8833 11583
rect 6897 11551 6903 11577
rect 6929 11551 6935 11577
rect 8807 11545 8833 11551
rect 9479 11577 9505 11583
rect 9479 11545 9505 11551
rect 10711 11577 10737 11583
rect 10711 11545 10737 11551
rect 11215 11577 11241 11583
rect 11887 11577 11913 11583
rect 11657 11551 11663 11577
rect 11689 11551 11695 11577
rect 12049 11551 12055 11577
rect 12081 11551 12087 11577
rect 12777 11551 12783 11577
rect 12809 11551 12815 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 11215 11545 11241 11551
rect 11887 11545 11913 11551
rect 8297 11495 8303 11521
rect 8329 11495 8335 11521
rect 10481 11495 10487 11521
rect 10513 11495 10519 11521
rect 13113 11495 13119 11521
rect 13145 11495 13151 11521
rect 14177 11495 14183 11521
rect 14209 11495 14215 11521
rect 11999 11465 12025 11471
rect 11999 11433 12025 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 10711 11297 10737 11303
rect 10711 11265 10737 11271
rect 12671 11297 12697 11303
rect 12671 11265 12697 11271
rect 13007 11297 13033 11303
rect 13007 11265 13033 11271
rect 10935 11241 10961 11247
rect 13399 11241 13425 11247
rect 11377 11215 11383 11241
rect 11409 11215 11415 11241
rect 11769 11215 11775 11241
rect 11801 11215 11807 11241
rect 10935 11209 10961 11215
rect 13399 11209 13425 11215
rect 8807 11185 8833 11191
rect 8807 11153 8833 11159
rect 9087 11185 9113 11191
rect 9087 11153 9113 11159
rect 9255 11185 9281 11191
rect 9255 11153 9281 11159
rect 9479 11185 9505 11191
rect 9479 11153 9505 11159
rect 9815 11185 9841 11191
rect 9815 11153 9841 11159
rect 10599 11185 10625 11191
rect 10599 11153 10625 11159
rect 12783 11185 12809 11191
rect 12783 11153 12809 11159
rect 12951 11185 12977 11191
rect 12951 11153 12977 11159
rect 13287 11185 13313 11191
rect 13287 11153 13313 11159
rect 13623 11185 13649 11191
rect 13623 11153 13649 11159
rect 13063 11129 13089 11135
rect 10033 11103 10039 11129
rect 10065 11103 10071 11129
rect 10313 11103 10319 11129
rect 10345 11103 10351 11129
rect 11489 11103 11495 11129
rect 11521 11103 11527 11129
rect 13063 11097 13089 11103
rect 13511 11129 13537 11135
rect 13511 11097 13537 11103
rect 13679 11129 13705 11135
rect 13679 11097 13705 11103
rect 13847 11129 13873 11135
rect 13847 11097 13873 11103
rect 13903 11129 13929 11135
rect 13903 11097 13929 11103
rect 14015 11129 14041 11135
rect 14015 11097 14041 11103
rect 8415 11073 8441 11079
rect 8415 11041 8441 11047
rect 9311 11073 9337 11079
rect 11999 11073 12025 11079
rect 12335 11073 12361 11079
rect 9865 11047 9871 11073
rect 9897 11047 9903 11073
rect 12161 11047 12167 11073
rect 12193 11047 12199 11073
rect 9311 11041 9337 11047
rect 11999 11041 12025 11047
rect 12335 11041 12361 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 6567 10905 6593 10911
rect 6567 10873 6593 10879
rect 8415 10905 8441 10911
rect 11657 10879 11663 10905
rect 11689 10879 11695 10905
rect 8415 10873 8441 10879
rect 8079 10849 8105 10855
rect 11831 10849 11857 10855
rect 8801 10823 8807 10849
rect 8833 10823 8839 10849
rect 14401 10823 14407 10849
rect 14433 10823 14439 10849
rect 8079 10817 8105 10823
rect 11831 10817 11857 10823
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 8297 10767 8303 10793
rect 8329 10767 8335 10793
rect 11321 10767 11327 10793
rect 11353 10767 11359 10793
rect 11545 10767 11551 10793
rect 11577 10767 11583 10793
rect 12049 10767 12055 10793
rect 12081 10767 12087 10793
rect 12609 10767 12615 10793
rect 12641 10767 12647 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 7961 10711 7967 10737
rect 7993 10711 7999 10737
rect 967 10681 993 10687
rect 967 10649 993 10655
rect 11887 10681 11913 10687
rect 20007 10681 20033 10687
rect 12329 10655 12335 10681
rect 12361 10655 12367 10681
rect 11887 10649 11913 10655
rect 20007 10649 20033 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 8577 10487 8583 10513
rect 8609 10487 8615 10513
rect 9143 10457 9169 10463
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 8185 10431 8191 10457
rect 8217 10431 8223 10457
rect 9143 10425 9169 10431
rect 9759 10457 9785 10463
rect 12609 10431 12615 10457
rect 12641 10431 12647 10457
rect 9759 10425 9785 10431
rect 9423 10401 9449 10407
rect 10151 10401 10177 10407
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 6785 10375 6791 10401
rect 6817 10375 6823 10401
rect 8577 10375 8583 10401
rect 8609 10375 8615 10401
rect 8801 10375 8807 10401
rect 8833 10375 8839 10401
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 9423 10369 9449 10375
rect 10151 10369 10177 10375
rect 10431 10401 10457 10407
rect 13679 10401 13705 10407
rect 10649 10375 10655 10401
rect 10681 10375 10687 10401
rect 10431 10369 10457 10375
rect 13679 10369 13705 10375
rect 13847 10401 13873 10407
rect 13847 10369 13873 10375
rect 13399 10345 13425 10351
rect 6057 10319 6063 10345
rect 6089 10319 6095 10345
rect 7121 10319 7127 10345
rect 7153 10319 7159 10345
rect 13399 10313 13425 10319
rect 13567 10345 13593 10351
rect 13567 10313 13593 10319
rect 13791 10345 13817 10351
rect 13791 10313 13817 10319
rect 9311 10289 9337 10295
rect 9311 10257 9337 10263
rect 9367 10289 9393 10295
rect 9367 10257 9393 10263
rect 9535 10289 9561 10295
rect 9535 10257 9561 10263
rect 13511 10289 13537 10295
rect 13511 10257 13537 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 6287 10121 6313 10127
rect 6287 10089 6313 10095
rect 7071 10121 7097 10127
rect 7071 10089 7097 10095
rect 14519 10121 14545 10127
rect 14519 10089 14545 10095
rect 6399 10065 6425 10071
rect 6399 10033 6425 10039
rect 6679 10065 6705 10071
rect 6679 10033 6705 10039
rect 7183 10065 7209 10071
rect 7183 10033 7209 10039
rect 7687 10065 7713 10071
rect 9143 10065 9169 10071
rect 8073 10039 8079 10065
rect 8105 10039 8111 10065
rect 8409 10039 8415 10065
rect 8441 10039 8447 10065
rect 9865 10039 9871 10065
rect 9897 10039 9903 10065
rect 10369 10039 10375 10065
rect 10401 10039 10407 10065
rect 12217 10039 12223 10065
rect 12249 10039 12255 10065
rect 13897 10039 13903 10065
rect 13929 10039 13935 10065
rect 7687 10033 7713 10039
rect 9143 10033 9169 10039
rect 6455 10009 6481 10015
rect 6455 9977 6481 9983
rect 6567 10009 6593 10015
rect 6567 9977 6593 9983
rect 6735 10009 6761 10015
rect 6735 9977 6761 9983
rect 7239 10009 7265 10015
rect 7239 9977 7265 9983
rect 7575 10009 7601 10015
rect 7575 9977 7601 9983
rect 7743 10009 7769 10015
rect 7743 9977 7769 9983
rect 7911 10009 7937 10015
rect 7911 9977 7937 9983
rect 8247 10009 8273 10015
rect 8247 9977 8273 9983
rect 8807 10009 8833 10015
rect 9255 10009 9281 10015
rect 12055 10009 12081 10015
rect 8969 9983 8975 10009
rect 9001 9983 9007 10009
rect 9585 9983 9591 10009
rect 9617 9983 9623 10009
rect 11209 9983 11215 10009
rect 11241 9983 11247 10009
rect 14289 9983 14295 10009
rect 14321 9983 14327 10009
rect 8807 9977 8833 9983
rect 9255 9977 9281 9983
rect 12055 9977 12081 9983
rect 10873 9927 10879 9953
rect 10905 9927 10911 9953
rect 12833 9927 12839 9953
rect 12865 9927 12871 9953
rect 9423 9897 9449 9903
rect 9423 9865 9449 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 10823 9729 10849 9735
rect 11433 9703 11439 9729
rect 11465 9703 11471 9729
rect 10823 9697 10849 9703
rect 9361 9647 9367 9673
rect 9393 9647 9399 9673
rect 9809 9647 9815 9673
rect 9841 9647 9847 9673
rect 10089 9647 10095 9673
rect 10121 9647 10127 9673
rect 10375 9617 10401 9623
rect 12111 9617 12137 9623
rect 8857 9591 8863 9617
rect 8889 9591 8895 9617
rect 9081 9591 9087 9617
rect 9113 9591 9119 9617
rect 9865 9591 9871 9617
rect 9897 9591 9903 9617
rect 11769 9591 11775 9617
rect 11801 9591 11807 9617
rect 10375 9585 10401 9591
rect 12111 9585 12137 9591
rect 12223 9617 12249 9623
rect 13231 9617 13257 9623
rect 12329 9591 12335 9617
rect 12361 9591 12367 9617
rect 13505 9591 13511 9617
rect 13537 9591 13543 9617
rect 12223 9585 12249 9591
rect 13231 9585 13257 9591
rect 10095 9561 10121 9567
rect 9137 9535 9143 9561
rect 9169 9535 9175 9561
rect 9753 9535 9759 9561
rect 9785 9535 9791 9561
rect 10095 9529 10121 9535
rect 10207 9561 10233 9567
rect 10207 9529 10233 9535
rect 10655 9561 10681 9567
rect 10655 9529 10681 9535
rect 10767 9561 10793 9567
rect 10767 9529 10793 9535
rect 13287 9505 13313 9511
rect 8745 9479 8751 9505
rect 8777 9479 8783 9505
rect 13287 9473 13313 9479
rect 13343 9505 13369 9511
rect 13343 9473 13369 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 14519 9337 14545 9343
rect 8241 9311 8247 9337
rect 8273 9311 8279 9337
rect 14519 9305 14545 9311
rect 7127 9281 7153 9287
rect 7127 9249 7153 9255
rect 7183 9281 7209 9287
rect 7183 9249 7209 9255
rect 11551 9281 11577 9287
rect 11551 9249 11577 9255
rect 7015 9225 7041 9231
rect 2137 9199 2143 9225
rect 2169 9199 2175 9225
rect 6897 9199 6903 9225
rect 6929 9199 6935 9225
rect 7015 9193 7041 9199
rect 8415 9225 8441 9231
rect 8415 9193 8441 9199
rect 8975 9225 9001 9231
rect 9871 9225 9897 9231
rect 9081 9199 9087 9225
rect 9113 9199 9119 9225
rect 8975 9193 9001 9199
rect 9871 9193 9897 9199
rect 10039 9225 10065 9231
rect 10039 9193 10065 9199
rect 10095 9225 10121 9231
rect 10095 9193 10121 9199
rect 10207 9225 10233 9231
rect 11383 9225 11409 9231
rect 11209 9199 11215 9225
rect 11241 9199 11247 9225
rect 10207 9193 10233 9199
rect 11383 9193 11409 9199
rect 11607 9225 11633 9231
rect 11607 9193 11633 9199
rect 11999 9225 12025 9231
rect 11999 9193 12025 9199
rect 12223 9225 12249 9231
rect 12223 9193 12249 9199
rect 12335 9225 12361 9231
rect 12335 9193 12361 9199
rect 12615 9225 12641 9231
rect 12833 9199 12839 9225
rect 12865 9199 12871 9225
rect 13225 9199 13231 9225
rect 13257 9199 13263 9225
rect 12615 9193 12641 9199
rect 7407 9169 7433 9175
rect 5441 9143 5447 9169
rect 5473 9143 5479 9169
rect 6505 9143 6511 9169
rect 6537 9143 6543 9169
rect 7407 9137 7433 9143
rect 9143 9169 9169 9175
rect 9143 9137 9169 9143
rect 11103 9169 11129 9175
rect 11103 9137 11129 9143
rect 11439 9169 11465 9175
rect 11439 9137 11465 9143
rect 12111 9169 12137 9175
rect 14289 9143 14295 9169
rect 14321 9143 14327 9169
rect 12111 9137 12137 9143
rect 967 9113 993 9119
rect 967 9081 993 9087
rect 11047 9113 11073 9119
rect 11047 9081 11073 9087
rect 12671 9113 12697 9119
rect 12671 9081 12697 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 10991 8945 11017 8951
rect 9641 8919 9647 8945
rect 9673 8919 9679 8945
rect 10991 8913 11017 8919
rect 967 8889 993 8895
rect 967 8857 993 8863
rect 10095 8889 10121 8895
rect 10095 8857 10121 8863
rect 10207 8889 10233 8895
rect 10207 8857 10233 8863
rect 11103 8889 11129 8895
rect 14631 8889 14657 8895
rect 14289 8863 14295 8889
rect 14321 8863 14327 8889
rect 11103 8857 11129 8863
rect 14631 8857 14657 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 6679 8833 6705 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6679 8801 6705 8807
rect 8023 8833 8049 8839
rect 9367 8833 9393 8839
rect 8241 8807 8247 8833
rect 8273 8807 8279 8833
rect 9081 8807 9087 8833
rect 9113 8807 9119 8833
rect 8023 8801 8049 8807
rect 9367 8801 9393 8807
rect 9535 8833 9561 8839
rect 11495 8833 11521 8839
rect 9753 8807 9759 8833
rect 9785 8807 9791 8833
rect 10761 8807 10767 8833
rect 10793 8807 10799 8833
rect 10873 8807 10879 8833
rect 10905 8807 10911 8833
rect 9535 8801 9561 8807
rect 11495 8801 11521 8807
rect 11607 8833 11633 8839
rect 11607 8801 11633 8807
rect 11663 8833 11689 8839
rect 11663 8801 11689 8807
rect 12055 8833 12081 8839
rect 12055 8801 12081 8807
rect 12391 8833 12417 8839
rect 12391 8801 12417 8807
rect 12503 8833 12529 8839
rect 12503 8801 12529 8807
rect 12727 8833 12753 8839
rect 12833 8807 12839 8833
rect 12865 8807 12871 8833
rect 18881 8807 18887 8833
rect 18913 8807 18919 8833
rect 12727 8801 12753 8807
rect 6791 8777 6817 8783
rect 6791 8745 6817 8751
rect 6847 8777 6873 8783
rect 6847 8745 6873 8751
rect 7239 8777 7265 8783
rect 7239 8745 7265 8751
rect 8079 8777 8105 8783
rect 8079 8745 8105 8751
rect 8135 8777 8161 8783
rect 8975 8777 9001 8783
rect 8297 8751 8303 8777
rect 8329 8751 8335 8777
rect 8135 8745 8161 8751
rect 8975 8745 9001 8751
rect 9199 8777 9225 8783
rect 9199 8745 9225 8751
rect 11215 8777 11241 8783
rect 11215 8745 11241 8751
rect 11383 8777 11409 8783
rect 12615 8777 12641 8783
rect 11881 8751 11887 8777
rect 11913 8751 11919 8777
rect 13225 8751 13231 8777
rect 13257 8751 13263 8777
rect 11383 8745 11409 8751
rect 12615 8745 12641 8751
rect 7295 8721 7321 8727
rect 7295 8689 7321 8695
rect 8919 8721 8945 8727
rect 8919 8689 8945 8695
rect 9423 8721 9449 8727
rect 11551 8721 11577 8727
rect 9921 8695 9927 8721
rect 9953 8695 9959 8721
rect 10929 8695 10935 8721
rect 10961 8695 10967 8721
rect 9423 8689 9449 8695
rect 11551 8689 11577 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 8919 8553 8945 8559
rect 8919 8521 8945 8527
rect 10991 8553 11017 8559
rect 10991 8521 11017 8527
rect 11327 8553 11353 8559
rect 11327 8521 11353 8527
rect 11663 8553 11689 8559
rect 11663 8521 11689 8527
rect 12055 8553 12081 8559
rect 12055 8521 12081 8527
rect 14463 8553 14489 8559
rect 14463 8521 14489 8527
rect 9031 8497 9057 8503
rect 7401 8471 7407 8497
rect 7433 8471 7439 8497
rect 9031 8465 9057 8471
rect 11439 8497 11465 8503
rect 11439 8465 11465 8471
rect 11943 8497 11969 8503
rect 11943 8465 11969 8471
rect 12167 8497 12193 8503
rect 13169 8471 13175 8497
rect 13201 8471 13207 8497
rect 12167 8465 12193 8471
rect 8023 8441 8049 8447
rect 8807 8441 8833 8447
rect 7793 8415 7799 8441
rect 7825 8415 7831 8441
rect 8689 8415 8695 8441
rect 8721 8415 8727 8441
rect 8023 8409 8049 8415
rect 8807 8409 8833 8415
rect 9255 8441 9281 8447
rect 9255 8409 9281 8415
rect 11103 8441 11129 8447
rect 12273 8415 12279 8441
rect 12305 8415 12311 8441
rect 12777 8415 12783 8441
rect 12809 8415 12815 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 11103 8409 11129 8415
rect 8863 8385 8889 8391
rect 6337 8359 6343 8385
rect 6369 8359 6375 8385
rect 8863 8353 8889 8359
rect 11719 8385 11745 8391
rect 11719 8353 11745 8359
rect 12111 8385 12137 8391
rect 20007 8385 20033 8391
rect 14233 8359 14239 8385
rect 14265 8359 14271 8385
rect 12111 8353 12137 8359
rect 20007 8353 20033 8359
rect 10935 8329 10961 8335
rect 10935 8297 10961 8303
rect 11271 8329 11297 8335
rect 11271 8297 11297 8303
rect 11775 8329 11801 8335
rect 11775 8297 11801 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 8807 8161 8833 8167
rect 8807 8129 8833 8135
rect 9199 8161 9225 8167
rect 9199 8129 9225 8135
rect 9311 8161 9337 8167
rect 9311 8129 9337 8135
rect 13847 8161 13873 8167
rect 13847 8129 13873 8135
rect 9647 8105 9673 8111
rect 14127 8105 14153 8111
rect 8633 8079 8639 8105
rect 8665 8079 8671 8105
rect 12553 8079 12559 8105
rect 12585 8079 12591 8105
rect 13617 8079 13623 8105
rect 13649 8079 13655 8105
rect 9647 8073 9673 8079
rect 14127 8073 14153 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 13791 8049 13817 8055
rect 7233 8023 7239 8049
rect 7265 8023 7271 8049
rect 8969 8023 8975 8049
rect 9001 8023 9007 8049
rect 9417 8023 9423 8049
rect 9449 8023 9455 8049
rect 9753 8023 9759 8049
rect 9785 8023 9791 8049
rect 12161 8023 12167 8049
rect 12193 8023 12199 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 13791 8017 13817 8023
rect 8863 7993 8889 7999
rect 7569 7967 7575 7993
rect 7601 7967 7607 7993
rect 8863 7961 8889 7967
rect 9143 7993 9169 7999
rect 9143 7961 9169 7967
rect 9591 7993 9617 7999
rect 9591 7961 9617 7967
rect 13847 7993 13873 7999
rect 13847 7961 13873 7967
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 13231 7769 13257 7775
rect 13231 7737 13257 7743
rect 13343 7769 13369 7775
rect 13343 7737 13369 7743
rect 13399 7713 13425 7719
rect 9081 7687 9087 7713
rect 9113 7687 9119 7713
rect 10817 7687 10823 7713
rect 10849 7687 10855 7713
rect 12049 7687 12055 7713
rect 12081 7687 12087 7713
rect 13399 7681 13425 7687
rect 12223 7657 12249 7663
rect 8745 7631 8751 7657
rect 8777 7631 8783 7657
rect 10481 7631 10487 7657
rect 10513 7631 10519 7657
rect 12223 7625 12249 7631
rect 10145 7575 10151 7601
rect 10177 7575 10183 7601
rect 11881 7575 11887 7601
rect 11913 7575 11919 7601
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 10319 7321 10345 7327
rect 10319 7289 10345 7295
rect 11999 7153 12025 7159
rect 11999 7121 12025 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 11775 6929 11801 6935
rect 11153 6903 11159 6929
rect 11185 6903 11191 6929
rect 11775 6897 11801 6903
rect 11489 6847 11495 6873
rect 11521 6847 11527 6873
rect 10089 6791 10095 6817
rect 10121 6791 10127 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 12391 2617 12417 2623
rect 12391 2585 12417 2591
rect 11881 2535 11887 2561
rect 11913 2535 11919 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9865 2143 9871 2169
rect 9897 2143 9903 2169
rect 10375 2057 10401 2063
rect 10375 2025 10401 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10705 1751 10711 1777
rect 10737 1751 10743 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 11215 1665 11241 1671
rect 11215 1633 11241 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 14687 19111 14713 19137
rect 9031 18999 9057 19025
rect 10711 18999 10737 19025
rect 12279 18999 12305 19025
rect 14295 18999 14321 19025
rect 8639 18943 8665 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 13119 18719 13145 18745
rect 14575 18719 14601 18745
rect 12615 18607 12641 18633
rect 14071 18607 14097 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 855 18159 881 18185
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 12223 14351 12249 14377
rect 10823 14295 10849 14321
rect 12391 14295 12417 14321
rect 11159 14239 11185 14265
rect 12559 14239 12585 14265
rect 12783 14239 12809 14265
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 11159 14015 11185 14041
rect 12279 14015 12305 14041
rect 2143 13903 2169 13929
rect 9311 13903 9337 13929
rect 11103 13903 11129 13929
rect 11215 13903 11241 13929
rect 11439 13903 11465 13929
rect 12167 13903 12193 13929
rect 12335 13903 12361 13929
rect 12615 13903 12641 13929
rect 9647 13847 9673 13873
rect 10711 13847 10737 13873
rect 10991 13847 11017 13873
rect 13007 13847 13033 13873
rect 14071 13847 14097 13873
rect 14295 13847 14321 13873
rect 967 13791 993 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 1023 13567 1049 13593
rect 12111 13567 12137 13593
rect 13791 13567 13817 13593
rect 2143 13511 2169 13537
rect 12055 13511 12081 13537
rect 12391 13511 12417 13537
rect 14015 13511 14041 13537
rect 7295 13455 7321 13481
rect 7463 13455 7489 13481
rect 9983 13455 10009 13481
rect 10151 13455 10177 13481
rect 12727 13455 12753 13481
rect 11943 13399 11969 13425
rect 12167 13399 12193 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7631 13231 7657 13257
rect 8919 13231 8945 13257
rect 9143 13231 9169 13257
rect 9255 13231 9281 13257
rect 10487 13231 10513 13257
rect 12671 13231 12697 13257
rect 12727 13231 12753 13257
rect 13119 13231 13145 13257
rect 13231 13231 13257 13257
rect 13511 13231 13537 13257
rect 13287 13175 13313 13201
rect 13567 13175 13593 13201
rect 2143 13119 2169 13145
rect 7407 13119 7433 13145
rect 7743 13119 7769 13145
rect 8695 13119 8721 13145
rect 8807 13119 8833 13145
rect 8975 13119 9001 13145
rect 9311 13119 9337 13145
rect 10431 13119 10457 13145
rect 10599 13119 10625 13145
rect 10711 13119 10737 13145
rect 12615 13119 12641 13145
rect 12951 13119 12977 13145
rect 13399 13119 13425 13145
rect 5951 13063 5977 13089
rect 7071 13063 7097 13089
rect 8023 13063 8049 13089
rect 8751 13063 8777 13089
rect 967 13007 993 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 6903 12839 6929 12865
rect 7967 12783 7993 12809
rect 9031 12783 9057 12809
rect 9255 12783 9281 12809
rect 11887 12783 11913 12809
rect 12167 12783 12193 12809
rect 20007 12783 20033 12809
rect 7631 12727 7657 12753
rect 10095 12727 10121 12753
rect 10207 12727 10233 12753
rect 10375 12727 10401 12753
rect 10935 12727 10961 12753
rect 11159 12727 11185 12753
rect 11663 12727 11689 12753
rect 11943 12727 11969 12753
rect 12055 12727 12081 12753
rect 12223 12727 12249 12753
rect 18831 12727 18857 12753
rect 6959 12671 6985 12697
rect 10655 12671 10681 12697
rect 11439 12671 11465 12697
rect 11775 12671 11801 12697
rect 12391 12671 12417 12697
rect 10711 12615 10737 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7239 12447 7265 12473
rect 7743 12447 7769 12473
rect 7799 12447 7825 12473
rect 8863 12447 8889 12473
rect 9143 12447 9169 12473
rect 11271 12447 11297 12473
rect 11663 12447 11689 12473
rect 12895 12447 12921 12473
rect 14911 12447 14937 12473
rect 7575 12391 7601 12417
rect 9871 12391 9897 12417
rect 7015 12335 7041 12361
rect 7687 12335 7713 12361
rect 7911 12335 7937 12361
rect 8695 12335 8721 12361
rect 9255 12335 9281 12361
rect 9479 12335 9505 12361
rect 11439 12335 11465 12361
rect 13063 12335 13089 12361
rect 13231 12335 13257 12361
rect 5559 12279 5585 12305
rect 6623 12279 6649 12305
rect 10935 12279 10961 12305
rect 13623 12279 13649 12305
rect 14687 12279 14713 12305
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 13847 12055 13873 12081
rect 967 11999 993 12025
rect 11271 11999 11297 12025
rect 11495 11999 11521 12025
rect 13399 11999 13425 12025
rect 2143 11943 2169 11969
rect 11159 11943 11185 11969
rect 13679 11943 13705 11969
rect 13791 11943 13817 11969
rect 6847 11887 6873 11913
rect 6903 11887 6929 11913
rect 7743 11887 7769 11913
rect 8191 11887 8217 11913
rect 13847 11887 13873 11913
rect 6735 11831 6761 11857
rect 7911 11831 7937 11857
rect 8023 11831 8049 11857
rect 8135 11831 8161 11857
rect 13343 11831 13369 11857
rect 13455 11831 13481 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 6511 11663 6537 11689
rect 6623 11663 6649 11689
rect 8639 11663 8665 11689
rect 8751 11663 8777 11689
rect 9311 11663 9337 11689
rect 14407 11663 14433 11689
rect 6679 11607 6705 11633
rect 7239 11607 7265 11633
rect 11047 11607 11073 11633
rect 11775 11607 11801 11633
rect 12167 11607 12193 11633
rect 6903 11551 6929 11577
rect 8807 11551 8833 11577
rect 9479 11551 9505 11577
rect 10711 11551 10737 11577
rect 11215 11551 11241 11577
rect 11663 11551 11689 11577
rect 11887 11551 11913 11577
rect 12055 11551 12081 11577
rect 12783 11551 12809 11577
rect 18831 11551 18857 11577
rect 8303 11495 8329 11521
rect 10487 11495 10513 11521
rect 13119 11495 13145 11521
rect 14183 11495 14209 11521
rect 11999 11439 12025 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 10711 11271 10737 11297
rect 12671 11271 12697 11297
rect 13007 11271 13033 11297
rect 10935 11215 10961 11241
rect 11383 11215 11409 11241
rect 11775 11215 11801 11241
rect 13399 11215 13425 11241
rect 8807 11159 8833 11185
rect 9087 11159 9113 11185
rect 9255 11159 9281 11185
rect 9479 11159 9505 11185
rect 9815 11159 9841 11185
rect 10599 11159 10625 11185
rect 12783 11159 12809 11185
rect 12951 11159 12977 11185
rect 13287 11159 13313 11185
rect 13623 11159 13649 11185
rect 10039 11103 10065 11129
rect 10319 11103 10345 11129
rect 11495 11103 11521 11129
rect 13063 11103 13089 11129
rect 13511 11103 13537 11129
rect 13679 11103 13705 11129
rect 13847 11103 13873 11129
rect 13903 11103 13929 11129
rect 14015 11103 14041 11129
rect 8415 11047 8441 11073
rect 9311 11047 9337 11073
rect 9871 11047 9897 11073
rect 11999 11047 12025 11073
rect 12167 11047 12193 11073
rect 12335 11047 12361 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 6567 10879 6593 10905
rect 8415 10879 8441 10905
rect 11663 10879 11689 10905
rect 8079 10823 8105 10849
rect 8807 10823 8833 10849
rect 11831 10823 11857 10849
rect 14407 10823 14433 10849
rect 2143 10767 2169 10793
rect 8303 10767 8329 10793
rect 11327 10767 11353 10793
rect 11551 10767 11577 10793
rect 12055 10767 12081 10793
rect 12615 10767 12641 10793
rect 18831 10767 18857 10793
rect 7967 10711 7993 10737
rect 967 10655 993 10681
rect 11887 10655 11913 10681
rect 12335 10655 12361 10681
rect 20007 10655 20033 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 8583 10487 8609 10513
rect 4999 10431 5025 10457
rect 8191 10431 8217 10457
rect 9143 10431 9169 10457
rect 9759 10431 9785 10457
rect 12615 10431 12641 10457
rect 6455 10375 6481 10401
rect 6791 10375 6817 10401
rect 8583 10375 8609 10401
rect 8807 10375 8833 10401
rect 9423 10375 9449 10401
rect 10039 10375 10065 10401
rect 10151 10375 10177 10401
rect 10431 10375 10457 10401
rect 10655 10375 10681 10401
rect 13679 10375 13705 10401
rect 13847 10375 13873 10401
rect 6063 10319 6089 10345
rect 7127 10319 7153 10345
rect 13399 10319 13425 10345
rect 13567 10319 13593 10345
rect 13791 10319 13817 10345
rect 9311 10263 9337 10289
rect 9367 10263 9393 10289
rect 9535 10263 9561 10289
rect 13511 10263 13537 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 6287 10095 6313 10121
rect 7071 10095 7097 10121
rect 14519 10095 14545 10121
rect 6399 10039 6425 10065
rect 6679 10039 6705 10065
rect 7183 10039 7209 10065
rect 7687 10039 7713 10065
rect 8079 10039 8105 10065
rect 8415 10039 8441 10065
rect 9143 10039 9169 10065
rect 9871 10039 9897 10065
rect 10375 10039 10401 10065
rect 12223 10039 12249 10065
rect 13903 10039 13929 10065
rect 6455 9983 6481 10009
rect 6567 9983 6593 10009
rect 6735 9983 6761 10009
rect 7239 9983 7265 10009
rect 7575 9983 7601 10009
rect 7743 9983 7769 10009
rect 7911 9983 7937 10009
rect 8247 9983 8273 10009
rect 8807 9983 8833 10009
rect 8975 9983 9001 10009
rect 9255 9983 9281 10009
rect 9591 9983 9617 10009
rect 11215 9983 11241 10009
rect 12055 9983 12081 10009
rect 14295 9983 14321 10009
rect 10879 9927 10905 9953
rect 12839 9927 12865 9953
rect 9423 9871 9449 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 10823 9703 10849 9729
rect 11439 9703 11465 9729
rect 9367 9647 9393 9673
rect 9815 9647 9841 9673
rect 10095 9647 10121 9673
rect 8863 9591 8889 9617
rect 9087 9591 9113 9617
rect 9871 9591 9897 9617
rect 10375 9591 10401 9617
rect 11775 9591 11801 9617
rect 12111 9591 12137 9617
rect 12223 9591 12249 9617
rect 12335 9591 12361 9617
rect 13231 9591 13257 9617
rect 13511 9591 13537 9617
rect 9143 9535 9169 9561
rect 9759 9535 9785 9561
rect 10095 9535 10121 9561
rect 10207 9535 10233 9561
rect 10655 9535 10681 9561
rect 10767 9535 10793 9561
rect 8751 9479 8777 9505
rect 13287 9479 13313 9505
rect 13343 9479 13369 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 8247 9311 8273 9337
rect 14519 9311 14545 9337
rect 7127 9255 7153 9281
rect 7183 9255 7209 9281
rect 11551 9255 11577 9281
rect 2143 9199 2169 9225
rect 6903 9199 6929 9225
rect 7015 9199 7041 9225
rect 8415 9199 8441 9225
rect 8975 9199 9001 9225
rect 9087 9199 9113 9225
rect 9871 9199 9897 9225
rect 10039 9199 10065 9225
rect 10095 9199 10121 9225
rect 10207 9199 10233 9225
rect 11215 9199 11241 9225
rect 11383 9199 11409 9225
rect 11607 9199 11633 9225
rect 11999 9199 12025 9225
rect 12223 9199 12249 9225
rect 12335 9199 12361 9225
rect 12615 9199 12641 9225
rect 12839 9199 12865 9225
rect 13231 9199 13257 9225
rect 5447 9143 5473 9169
rect 6511 9143 6537 9169
rect 7407 9143 7433 9169
rect 9143 9143 9169 9169
rect 11103 9143 11129 9169
rect 11439 9143 11465 9169
rect 12111 9143 12137 9169
rect 14295 9143 14321 9169
rect 967 9087 993 9113
rect 11047 9087 11073 9113
rect 12671 9087 12697 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 9647 8919 9673 8945
rect 10991 8919 11017 8945
rect 967 8863 993 8889
rect 10095 8863 10121 8889
rect 10207 8863 10233 8889
rect 11103 8863 11129 8889
rect 14295 8863 14321 8889
rect 14631 8863 14657 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 6679 8807 6705 8833
rect 8023 8807 8049 8833
rect 8247 8807 8273 8833
rect 9087 8807 9113 8833
rect 9367 8807 9393 8833
rect 9535 8807 9561 8833
rect 9759 8807 9785 8833
rect 10767 8807 10793 8833
rect 10879 8807 10905 8833
rect 11495 8807 11521 8833
rect 11607 8807 11633 8833
rect 11663 8807 11689 8833
rect 12055 8807 12081 8833
rect 12391 8807 12417 8833
rect 12503 8807 12529 8833
rect 12727 8807 12753 8833
rect 12839 8807 12865 8833
rect 18887 8807 18913 8833
rect 6791 8751 6817 8777
rect 6847 8751 6873 8777
rect 7239 8751 7265 8777
rect 8079 8751 8105 8777
rect 8135 8751 8161 8777
rect 8303 8751 8329 8777
rect 8975 8751 9001 8777
rect 9199 8751 9225 8777
rect 11215 8751 11241 8777
rect 11383 8751 11409 8777
rect 11887 8751 11913 8777
rect 12615 8751 12641 8777
rect 13231 8751 13257 8777
rect 7295 8695 7321 8721
rect 8919 8695 8945 8721
rect 9423 8695 9449 8721
rect 9927 8695 9953 8721
rect 10935 8695 10961 8721
rect 11551 8695 11577 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 8919 8527 8945 8553
rect 10991 8527 11017 8553
rect 11327 8527 11353 8553
rect 11663 8527 11689 8553
rect 12055 8527 12081 8553
rect 14463 8527 14489 8553
rect 7407 8471 7433 8497
rect 9031 8471 9057 8497
rect 11439 8471 11465 8497
rect 11943 8471 11969 8497
rect 12167 8471 12193 8497
rect 13175 8471 13201 8497
rect 7799 8415 7825 8441
rect 8023 8415 8049 8441
rect 8695 8415 8721 8441
rect 8807 8415 8833 8441
rect 9255 8415 9281 8441
rect 11103 8415 11129 8441
rect 12279 8415 12305 8441
rect 12783 8415 12809 8441
rect 18831 8415 18857 8441
rect 6343 8359 6369 8385
rect 8863 8359 8889 8385
rect 11719 8359 11745 8385
rect 12111 8359 12137 8385
rect 14239 8359 14265 8385
rect 20007 8359 20033 8385
rect 10935 8303 10961 8329
rect 11271 8303 11297 8329
rect 11775 8303 11801 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 8807 8135 8833 8161
rect 9199 8135 9225 8161
rect 9311 8135 9337 8161
rect 13847 8135 13873 8161
rect 8639 8079 8665 8105
rect 9647 8079 9673 8105
rect 12559 8079 12585 8105
rect 13623 8079 13649 8105
rect 14127 8079 14153 8105
rect 20007 8079 20033 8105
rect 7239 8023 7265 8049
rect 8975 8023 9001 8049
rect 9423 8023 9449 8049
rect 9759 8023 9785 8049
rect 12167 8023 12193 8049
rect 13791 8023 13817 8049
rect 18831 8023 18857 8049
rect 7575 7967 7601 7993
rect 8863 7967 8889 7993
rect 9143 7967 9169 7993
rect 9591 7967 9617 7993
rect 13847 7967 13873 7993
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 13231 7743 13257 7769
rect 13343 7743 13369 7769
rect 9087 7687 9113 7713
rect 10823 7687 10849 7713
rect 12055 7687 12081 7713
rect 13399 7687 13425 7713
rect 8751 7631 8777 7657
rect 10487 7631 10513 7657
rect 12223 7631 12249 7657
rect 10151 7575 10177 7601
rect 11887 7575 11913 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 10319 7295 10345 7321
rect 11999 7127 12025 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 11159 6903 11185 6929
rect 11775 6903 11801 6929
rect 11495 6847 11521 6873
rect 10095 6791 10121 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 12391 2591 12417 2617
rect 11887 2535 11913 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9871 2143 9897 2169
rect 10375 2031 10401 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 12783 1807 12809 1833
rect 8807 1751 8833 1777
rect 10711 1751 10737 1777
rect 12279 1751 12305 1777
rect 11215 1639 11241 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8736 20600 8792 21000
rect 9072 20600 9128 21000
rect 10752 20600 10808 21000
rect 12096 20600 12152 21000
rect 12432 20600 12488 21000
rect 13440 20600 13496 21000
rect 13776 20600 13832 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8638 18970 8666 18975
rect 8750 18970 8778 20600
rect 9086 19138 9114 20600
rect 9310 19138 9338 19143
rect 9086 19137 9338 19138
rect 9086 19111 9311 19137
rect 9337 19111 9338 19137
rect 9086 19110 9338 19111
rect 9310 19105 9338 19110
rect 10766 19138 10794 20600
rect 10766 19105 10794 19110
rect 11214 19138 11242 19143
rect 11214 19091 11242 19110
rect 12110 19138 12138 20600
rect 12110 19105 12138 19110
rect 8638 18969 8778 18970
rect 8638 18943 8639 18969
rect 8665 18943 8778 18969
rect 8638 18942 8778 18943
rect 9030 19025 9058 19031
rect 9030 18999 9031 19025
rect 9057 18999 9058 19025
rect 8638 18937 8666 18942
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 854 18186 882 18191
rect 854 18139 882 18158
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 9030 15974 9058 18999
rect 10710 19025 10738 19031
rect 10710 18999 10711 19025
rect 10737 18999 10738 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9030 15946 9226 15974
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2086 14154 2114 14159
rect 966 13817 994 13823
rect 966 13791 967 13817
rect 993 13791 994 13817
rect 966 13482 994 13791
rect 966 13449 994 13454
rect 1022 13593 1050 13599
rect 1022 13567 1023 13593
rect 1049 13567 1050 13593
rect 1022 13146 1050 13567
rect 1022 13113 1050 13118
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 10681 994 10687
rect 966 10655 967 10681
rect 993 10655 994 10681
rect 966 10458 994 10655
rect 966 10425 994 10430
rect 2086 10290 2114 14126
rect 2142 13930 2170 13935
rect 2142 13883 2170 13902
rect 7630 13930 7658 13935
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 2142 13538 2170 13543
rect 2142 13491 2170 13510
rect 7294 13538 7322 13543
rect 7294 13481 7322 13510
rect 7294 13455 7295 13481
rect 7321 13455 7322 13481
rect 7294 13449 7322 13455
rect 7462 13481 7490 13487
rect 7462 13455 7463 13481
rect 7489 13455 7490 13481
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 5950 13146 5978 13151
rect 5950 13089 5978 13118
rect 7406 13145 7434 13151
rect 7406 13119 7407 13145
rect 7433 13119 7434 13145
rect 7070 13090 7098 13095
rect 7406 13090 7434 13119
rect 7462 13146 7490 13455
rect 7630 13257 7658 13902
rect 8918 13818 8946 13823
rect 7630 13231 7631 13257
rect 7657 13231 7658 13257
rect 7630 13225 7658 13231
rect 8862 13790 8918 13818
rect 7742 13146 7770 13151
rect 7490 13118 7602 13146
rect 7462 13113 7490 13118
rect 5950 13063 5951 13089
rect 5977 13063 5978 13089
rect 5950 13057 5978 13063
rect 6902 13089 7098 13090
rect 6902 13063 7071 13089
rect 7097 13063 7098 13089
rect 6902 13062 7098 13063
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6902 12865 6930 13062
rect 7070 13057 7098 13062
rect 7238 13062 7406 13090
rect 6902 12839 6903 12865
rect 6929 12839 6930 12865
rect 6902 12833 6930 12839
rect 6958 12697 6986 12703
rect 6958 12671 6959 12697
rect 6985 12671 6986 12697
rect 6958 12474 6986 12671
rect 7238 12474 7266 13062
rect 7406 13057 7434 13062
rect 6958 12441 6986 12446
rect 7014 12473 7266 12474
rect 7014 12447 7239 12473
rect 7265 12447 7266 12473
rect 7014 12446 7266 12447
rect 7014 12362 7042 12446
rect 7238 12441 7266 12446
rect 7574 12417 7602 13118
rect 7742 13099 7770 13118
rect 8694 13146 8722 13151
rect 8694 13099 8722 13118
rect 8806 13145 8834 13151
rect 8806 13119 8807 13145
rect 8833 13119 8834 13145
rect 7630 13090 7658 13095
rect 7630 12753 7658 13062
rect 8022 13090 8050 13095
rect 8022 13043 8050 13062
rect 8750 13089 8778 13095
rect 8750 13063 8751 13089
rect 8777 13063 8778 13089
rect 7966 12810 7994 12815
rect 7966 12763 7994 12782
rect 8750 12810 8778 13063
rect 8750 12777 8778 12782
rect 7630 12727 7631 12753
rect 7657 12727 7658 12753
rect 7630 12721 7658 12727
rect 7798 12530 7826 12535
rect 7742 12474 7770 12479
rect 7742 12427 7770 12446
rect 7798 12473 7826 12502
rect 8806 12530 8834 13119
rect 8862 13146 8890 13790
rect 8918 13785 8946 13790
rect 8918 13258 8946 13263
rect 9142 13258 9170 13263
rect 8918 13257 9170 13258
rect 8918 13231 8919 13257
rect 8945 13231 9143 13257
rect 9169 13231 9170 13257
rect 8918 13230 9170 13231
rect 8918 13225 8946 13230
rect 9142 13225 9170 13230
rect 9198 13258 9226 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9310 13930 9338 13935
rect 10654 13930 10682 13935
rect 9310 13929 9394 13930
rect 9310 13903 9311 13929
rect 9337 13903 9394 13929
rect 9310 13902 9394 13903
rect 9310 13897 9338 13902
rect 9366 13874 9394 13902
rect 9254 13258 9282 13263
rect 9198 13257 9282 13258
rect 9198 13231 9255 13257
rect 9281 13231 9282 13257
rect 9198 13230 9282 13231
rect 8974 13146 9002 13151
rect 9142 13146 9170 13151
rect 8862 13145 9002 13146
rect 8862 13119 8975 13145
rect 9001 13119 9002 13145
rect 8862 13118 9002 13119
rect 8806 12497 8834 12502
rect 7798 12447 7799 12473
rect 7825 12447 7826 12473
rect 7798 12441 7826 12447
rect 7910 12474 7938 12479
rect 7574 12391 7575 12417
rect 7601 12391 7602 12417
rect 7574 12385 7602 12391
rect 6958 12361 7042 12362
rect 6958 12335 7015 12361
rect 7041 12335 7042 12361
rect 6958 12334 7042 12335
rect 5558 12305 5586 12311
rect 6622 12306 6650 12311
rect 5558 12279 5559 12305
rect 5585 12279 5586 12305
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 5558 11970 5586 12279
rect 5558 11937 5586 11942
rect 6510 12305 6650 12306
rect 6510 12279 6623 12305
rect 6649 12279 6650 12305
rect 6510 12278 6650 12279
rect 6510 11689 6538 12278
rect 6622 12273 6650 12278
rect 6846 11970 6874 11975
rect 6846 11913 6874 11942
rect 6846 11887 6847 11913
rect 6873 11887 6874 11913
rect 6846 11881 6874 11887
rect 6902 11914 6930 11919
rect 6734 11858 6762 11863
rect 6678 11857 6762 11858
rect 6678 11831 6735 11857
rect 6761 11831 6762 11857
rect 6678 11830 6762 11831
rect 6510 11663 6511 11689
rect 6537 11663 6538 11689
rect 6510 11657 6538 11663
rect 6622 11690 6650 11695
rect 6622 11643 6650 11662
rect 6678 11633 6706 11830
rect 6734 11825 6762 11830
rect 6902 11690 6930 11886
rect 6678 11607 6679 11633
rect 6705 11607 6706 11633
rect 6678 11601 6706 11607
rect 6846 11662 6930 11690
rect 6846 11578 6874 11662
rect 6734 11550 6874 11578
rect 6902 11578 6930 11583
rect 6958 11578 6986 12334
rect 7014 12329 7042 12334
rect 7686 12362 7714 12367
rect 7686 12361 7770 12362
rect 7686 12335 7687 12361
rect 7713 12335 7770 12361
rect 7686 12334 7770 12335
rect 7686 12329 7714 12334
rect 7742 11914 7770 12334
rect 7910 12361 7938 12446
rect 8862 12474 8890 12479
rect 8918 12474 8946 13118
rect 8974 13113 9002 13118
rect 9086 13118 9142 13146
rect 9030 13034 9058 13039
rect 9030 12809 9058 13006
rect 9030 12783 9031 12809
rect 9057 12783 9058 12809
rect 9030 12777 9058 12783
rect 8862 12473 8946 12474
rect 8862 12447 8863 12473
rect 8889 12447 8946 12473
rect 8862 12446 8946 12447
rect 9086 12474 9114 13118
rect 9142 13113 9170 13118
rect 9198 13034 9226 13230
rect 9254 13225 9282 13230
rect 9198 13001 9226 13006
rect 9310 13145 9338 13151
rect 9310 13119 9311 13145
rect 9337 13119 9338 13145
rect 9310 13034 9338 13119
rect 9310 13001 9338 13006
rect 9366 13090 9394 13846
rect 9646 13874 9674 13879
rect 9646 13873 10010 13874
rect 9646 13847 9647 13873
rect 9673 13847 10010 13873
rect 9646 13846 10010 13847
rect 9646 13841 9674 13846
rect 9982 13481 10010 13846
rect 9982 13455 9983 13481
rect 10009 13455 10010 13481
rect 9982 13449 10010 13455
rect 10150 13481 10178 13487
rect 10150 13455 10151 13481
rect 10177 13455 10178 13481
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9366 12866 9394 13062
rect 9534 13034 9562 13039
rect 9254 12838 9506 12866
rect 9254 12809 9282 12838
rect 9254 12783 9255 12809
rect 9281 12783 9282 12809
rect 9254 12777 9282 12783
rect 9142 12474 9170 12479
rect 9114 12473 9170 12474
rect 9114 12447 9143 12473
rect 9169 12447 9170 12473
rect 9114 12446 9170 12447
rect 8862 12441 8890 12446
rect 9086 12427 9114 12446
rect 9142 12441 9170 12446
rect 8694 12362 8722 12367
rect 7910 12335 7911 12361
rect 7937 12335 7938 12361
rect 7910 12329 7938 12335
rect 8526 12361 8722 12362
rect 8526 12335 8695 12361
rect 8721 12335 8722 12361
rect 8526 12334 8722 12335
rect 7742 11867 7770 11886
rect 8190 11913 8218 11919
rect 8190 11887 8191 11913
rect 8217 11887 8218 11913
rect 7238 11858 7266 11863
rect 7238 11633 7266 11830
rect 7238 11607 7239 11633
rect 7265 11607 7266 11633
rect 7238 11601 7266 11607
rect 7910 11857 7938 11863
rect 7910 11831 7911 11857
rect 7937 11831 7938 11857
rect 6902 11577 6986 11578
rect 6902 11551 6903 11577
rect 6929 11551 6986 11577
rect 6902 11550 6986 11551
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 6566 10906 6594 10911
rect 6454 10878 6566 10906
rect 2142 10794 2170 10799
rect 2142 10747 2170 10766
rect 4998 10794 5026 10799
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 4998 10458 5026 10766
rect 4998 10411 5026 10430
rect 6454 10401 6482 10878
rect 6566 10859 6594 10878
rect 6454 10375 6455 10401
rect 6481 10375 6482 10401
rect 6454 10369 6482 10375
rect 6678 10458 6706 10463
rect 6062 10346 6090 10351
rect 6062 10345 6314 10346
rect 6062 10319 6063 10345
rect 6089 10319 6314 10345
rect 6062 10318 6314 10319
rect 6062 10313 6090 10318
rect 2086 10257 2114 10262
rect 6286 10121 6314 10318
rect 6286 10095 6287 10121
rect 6313 10095 6314 10121
rect 6286 10089 6314 10095
rect 6398 10066 6426 10071
rect 6398 10019 6426 10038
rect 6678 10065 6706 10430
rect 6678 10039 6679 10065
rect 6705 10039 6706 10065
rect 6678 10033 6706 10039
rect 6454 10010 6482 10015
rect 6566 10010 6594 10015
rect 6454 10009 6594 10010
rect 6454 9983 6455 10009
rect 6481 9983 6567 10009
rect 6593 9983 6594 10009
rect 6454 9982 6594 9983
rect 6454 9977 6482 9982
rect 6566 9977 6594 9982
rect 6734 10009 6762 11550
rect 6902 10906 6930 11550
rect 6790 10878 6902 10906
rect 6790 10401 6818 10878
rect 6902 10873 6930 10878
rect 7910 10514 7938 11831
rect 8022 11858 8050 11863
rect 8022 11811 8050 11830
rect 8134 11857 8162 11863
rect 8134 11831 8135 11857
rect 8161 11831 8162 11857
rect 8078 11690 8106 11695
rect 8134 11690 8162 11831
rect 8106 11662 8162 11690
rect 8190 11690 8218 11887
rect 8078 11657 8106 11662
rect 8190 11657 8218 11662
rect 8302 11521 8330 11527
rect 8302 11495 8303 11521
rect 8329 11495 8330 11521
rect 8302 11186 8330 11495
rect 8302 11130 8330 11158
rect 8190 11102 8330 11130
rect 8078 10850 8106 10855
rect 8190 10850 8218 11102
rect 8414 11074 8442 11079
rect 8414 11073 8498 11074
rect 8414 11047 8415 11073
rect 8441 11047 8498 11073
rect 8414 11046 8498 11047
rect 8414 11041 8442 11046
rect 8414 10906 8442 10911
rect 8414 10859 8442 10878
rect 8078 10849 8218 10850
rect 8078 10823 8079 10849
rect 8105 10823 8218 10849
rect 8078 10822 8218 10823
rect 8470 10850 8498 11046
rect 8078 10817 8106 10822
rect 8470 10817 8498 10822
rect 8302 10794 8330 10799
rect 8302 10747 8330 10766
rect 7910 10481 7938 10486
rect 7966 10737 7994 10743
rect 7966 10711 7967 10737
rect 7993 10711 7994 10737
rect 6790 10375 6791 10401
rect 6817 10375 6818 10401
rect 6790 10094 6818 10375
rect 7966 10402 7994 10711
rect 7126 10346 7154 10351
rect 7070 10345 7154 10346
rect 7070 10319 7127 10345
rect 7153 10319 7154 10345
rect 7070 10318 7154 10319
rect 7070 10121 7098 10318
rect 7126 10313 7154 10318
rect 7798 10234 7826 10239
rect 7070 10095 7071 10121
rect 7097 10095 7098 10121
rect 6790 10066 6930 10094
rect 7070 10089 7098 10095
rect 7742 10122 7770 10127
rect 6734 9983 6735 10009
rect 6761 9983 6762 10009
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 6734 9282 6762 9983
rect 6734 9249 6762 9254
rect 2142 9226 2170 9231
rect 2142 9179 2170 9198
rect 5446 9226 5474 9231
rect 5446 9169 5474 9198
rect 6902 9225 6930 10066
rect 7182 10066 7210 10071
rect 7182 9786 7210 10038
rect 7686 10066 7770 10094
rect 7686 10065 7714 10066
rect 7686 10039 7687 10065
rect 7713 10039 7714 10065
rect 7686 10033 7714 10039
rect 7238 10010 7266 10015
rect 7238 9963 7266 9982
rect 7574 10010 7602 10015
rect 7574 9963 7602 9982
rect 7742 10010 7770 10015
rect 7798 10010 7826 10206
rect 7742 10009 7826 10010
rect 7742 9983 7743 10009
rect 7769 9983 7826 10009
rect 7742 9982 7826 9983
rect 7910 10010 7938 10015
rect 7742 9977 7770 9982
rect 7910 9963 7938 9982
rect 7182 9753 7210 9758
rect 7126 9281 7154 9287
rect 7126 9255 7127 9281
rect 7153 9255 7154 9281
rect 7014 9226 7042 9231
rect 6902 9199 6903 9225
rect 6929 9199 6930 9225
rect 5446 9143 5447 9169
rect 5473 9143 5474 9169
rect 5446 9137 5474 9143
rect 6510 9170 6538 9175
rect 6902 9170 6930 9199
rect 6510 9169 6706 9170
rect 6510 9143 6511 9169
rect 6537 9143 6706 9169
rect 6510 9142 6706 9143
rect 6510 9137 6538 9142
rect 966 9114 994 9119
rect 966 9067 994 9086
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8889 994 8895
rect 966 8863 967 8889
rect 993 8863 994 8889
rect 966 8442 994 8863
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 6342 8834 6370 8839
rect 966 8409 994 8414
rect 6342 8385 6370 8806
rect 6678 8833 6706 9142
rect 6902 9137 6930 9142
rect 6958 9225 7042 9226
rect 6958 9199 7015 9225
rect 7041 9199 7042 9225
rect 6958 9198 7042 9199
rect 6958 8890 6986 9198
rect 7014 9193 7042 9198
rect 7126 9226 7154 9255
rect 7182 9282 7210 9287
rect 7182 9235 7210 9254
rect 7126 9193 7154 9198
rect 7406 9170 7434 9175
rect 7434 9142 7490 9170
rect 7406 9123 7434 9142
rect 6678 8807 6679 8833
rect 6705 8807 6706 8833
rect 6678 8801 6706 8807
rect 6790 8862 6986 8890
rect 6790 8777 6818 8862
rect 6790 8751 6791 8777
rect 6817 8751 6818 8777
rect 6790 8745 6818 8751
rect 6846 8777 6874 8783
rect 6846 8751 6847 8777
rect 6873 8751 6874 8777
rect 6846 8722 6874 8751
rect 7238 8778 7266 8783
rect 7238 8731 7266 8750
rect 6846 8689 6874 8694
rect 7294 8722 7322 8727
rect 7294 8721 7434 8722
rect 7294 8695 7295 8721
rect 7321 8695 7434 8721
rect 7294 8694 7434 8695
rect 7294 8689 7322 8694
rect 7406 8497 7434 8694
rect 7406 8471 7407 8497
rect 7433 8471 7434 8497
rect 7406 8465 7434 8471
rect 6342 8359 6343 8385
rect 6369 8359 6370 8385
rect 6342 8353 6370 8359
rect 7238 8442 7266 8447
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 7238 8049 7266 8414
rect 7462 8442 7490 9142
rect 7966 8834 7994 10374
rect 8190 10457 8218 10463
rect 8190 10431 8191 10457
rect 8217 10431 8218 10457
rect 8078 10066 8106 10071
rect 8078 10019 8106 10038
rect 8190 10010 8218 10431
rect 8526 10178 8554 12334
rect 8694 12329 8722 12334
rect 9254 12361 9282 12367
rect 9254 12335 9255 12361
rect 9281 12335 9282 12361
rect 8638 11690 8666 11695
rect 8638 11643 8666 11662
rect 8750 11690 8778 11695
rect 8750 11643 8778 11662
rect 8806 11578 8834 11583
rect 8694 11577 8834 11578
rect 8694 11551 8807 11577
rect 8833 11551 8834 11577
rect 8694 11550 8834 11551
rect 8582 10514 8610 10519
rect 8582 10467 8610 10486
rect 8582 10402 8610 10407
rect 8582 10355 8610 10374
rect 8694 10234 8722 11550
rect 8806 11545 8834 11550
rect 9254 11298 9282 12335
rect 9478 12361 9506 12838
rect 9478 12335 9479 12361
rect 9505 12335 9506 12361
rect 9478 12329 9506 12335
rect 9534 12250 9562 13006
rect 10094 12753 10122 12759
rect 10094 12727 10095 12753
rect 10121 12727 10122 12753
rect 9918 12558 10050 12563
rect 9646 12530 9674 12535
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9674 12502 9730 12530
rect 9918 12525 10050 12530
rect 9646 12497 9674 12502
rect 9310 12222 9562 12250
rect 9310 11690 9338 12222
rect 9310 11643 9338 11662
rect 9478 11578 9506 11583
rect 9478 11577 9618 11578
rect 9478 11551 9479 11577
rect 9505 11551 9618 11577
rect 9478 11550 9618 11551
rect 9478 11545 9506 11550
rect 9254 11270 9338 11298
rect 8806 11186 8834 11191
rect 8694 10201 8722 10206
rect 8750 11185 8834 11186
rect 8750 11159 8807 11185
rect 8833 11159 8834 11185
rect 8750 11158 8834 11159
rect 8750 10794 8778 11158
rect 8806 11153 8834 11158
rect 9086 11186 9114 11191
rect 9254 11186 9282 11191
rect 9114 11185 9282 11186
rect 9114 11159 9255 11185
rect 9281 11159 9282 11185
rect 9114 11158 9282 11159
rect 9086 11139 9114 11158
rect 9254 11153 9282 11158
rect 9310 11186 9338 11270
rect 9310 11073 9338 11158
rect 9310 11047 9311 11073
rect 9337 11047 9338 11073
rect 9310 11041 9338 11047
rect 9478 11185 9506 11191
rect 9478 11159 9479 11185
rect 9505 11159 9506 11185
rect 9422 10962 9450 10967
rect 8806 10850 8834 10855
rect 8806 10803 8834 10822
rect 9142 10850 9170 10855
rect 8246 10150 8554 10178
rect 8246 10122 8274 10150
rect 8750 10122 8778 10766
rect 9142 10458 9170 10822
rect 9142 10457 9226 10458
rect 9142 10431 9143 10457
rect 9169 10431 9226 10457
rect 9142 10430 9226 10431
rect 9142 10425 9170 10430
rect 8806 10402 8834 10407
rect 9086 10402 9114 10407
rect 8806 10401 8946 10402
rect 8806 10375 8807 10401
rect 8833 10375 8946 10401
rect 8806 10374 8946 10375
rect 8806 10369 8834 10374
rect 8246 10066 8330 10094
rect 8750 10089 8778 10094
rect 8918 10094 8946 10374
rect 8190 9977 8218 9982
rect 8246 10009 8274 10015
rect 8246 9983 8247 10009
rect 8273 9983 8274 10009
rect 8246 9954 8274 9983
rect 8246 9921 8274 9926
rect 8246 9338 8274 9343
rect 8302 9338 8330 10066
rect 8246 9337 8330 9338
rect 8246 9311 8247 9337
rect 8273 9311 8330 9337
rect 8246 9310 8330 9311
rect 8246 9305 8274 9310
rect 8022 8834 8050 8839
rect 7966 8833 8050 8834
rect 7966 8807 8023 8833
rect 8049 8807 8050 8833
rect 7966 8806 8050 8807
rect 8022 8801 8050 8806
rect 8134 8834 8162 8839
rect 8078 8778 8106 8783
rect 8078 8731 8106 8750
rect 8134 8777 8162 8806
rect 8246 8834 8274 8839
rect 8246 8787 8274 8806
rect 8134 8751 8135 8777
rect 8161 8751 8162 8777
rect 8134 8745 8162 8751
rect 8302 8778 8330 9310
rect 8414 10065 8442 10071
rect 8414 10039 8415 10065
rect 8441 10039 8442 10065
rect 8414 9338 8442 10039
rect 8862 10066 8890 10071
rect 8918 10066 9002 10094
rect 8806 10010 8834 10015
rect 8806 9963 8834 9982
rect 8862 9617 8890 10038
rect 8974 10010 9002 10066
rect 8974 9963 9002 9982
rect 8862 9591 8863 9617
rect 8889 9591 8890 9617
rect 8862 9585 8890 9591
rect 9086 9617 9114 10374
rect 9086 9591 9087 9617
rect 9113 9591 9114 9617
rect 8414 9305 8442 9310
rect 8750 9505 8778 9511
rect 8750 9479 8751 9505
rect 8777 9479 8778 9505
rect 8414 9226 8442 9231
rect 8414 9179 8442 9198
rect 8750 9226 8778 9479
rect 8750 9193 8778 9198
rect 8918 9338 8946 9343
rect 8918 9114 8946 9310
rect 8974 9226 9002 9231
rect 8974 9179 9002 9198
rect 9086 9225 9114 9591
rect 9142 10066 9170 10071
rect 9142 9898 9170 10038
rect 9198 9898 9226 10430
rect 9422 10401 9450 10934
rect 9422 10375 9423 10401
rect 9449 10375 9450 10401
rect 9422 10369 9450 10375
rect 9310 10346 9338 10351
rect 9310 10289 9338 10318
rect 9310 10263 9311 10289
rect 9337 10263 9338 10289
rect 9310 10234 9338 10263
rect 9310 10201 9338 10206
rect 9366 10289 9394 10295
rect 9366 10263 9367 10289
rect 9393 10263 9394 10289
rect 9254 10122 9282 10127
rect 9254 10009 9282 10094
rect 9366 10066 9394 10263
rect 9254 9983 9255 10009
rect 9281 9983 9282 10009
rect 9254 9977 9282 9983
rect 9310 10038 9394 10066
rect 9198 9870 9282 9898
rect 9142 9561 9170 9870
rect 9142 9535 9143 9561
rect 9169 9535 9170 9561
rect 9142 9529 9170 9535
rect 9198 9562 9226 9567
rect 9086 9199 9087 9225
rect 9113 9199 9114 9225
rect 9086 9193 9114 9199
rect 9142 9169 9170 9175
rect 9142 9143 9143 9169
rect 9169 9143 9170 9169
rect 9142 9114 9170 9143
rect 8918 9086 9002 9114
rect 8302 8731 8330 8750
rect 8694 8778 8722 8783
rect 7462 8409 7490 8414
rect 7798 8442 7826 8447
rect 7798 8395 7826 8414
rect 8022 8442 8050 8447
rect 8022 8395 8050 8414
rect 8694 8441 8722 8750
rect 8974 8777 9002 9086
rect 8974 8751 8975 8777
rect 9001 8751 9002 8777
rect 8974 8745 9002 8751
rect 9030 9086 9142 9114
rect 8918 8722 8946 8727
rect 8918 8675 8946 8694
rect 9030 8610 9058 9086
rect 9142 9081 9170 9086
rect 9198 9002 9226 9534
rect 9086 8974 9226 9002
rect 9086 8833 9114 8974
rect 9086 8807 9087 8833
rect 9113 8807 9114 8833
rect 9086 8801 9114 8807
rect 9198 8834 9226 8839
rect 8918 8582 9058 8610
rect 9142 8778 9170 8783
rect 8918 8553 8946 8582
rect 8918 8527 8919 8553
rect 8945 8527 8946 8553
rect 8918 8521 8946 8527
rect 9030 8498 9058 8503
rect 9142 8498 9170 8750
rect 9198 8777 9226 8806
rect 9198 8751 9199 8777
rect 9225 8751 9226 8777
rect 9198 8722 9226 8751
rect 9198 8689 9226 8694
rect 9030 8497 9170 8498
rect 9030 8471 9031 8497
rect 9057 8471 9170 8497
rect 9030 8470 9170 8471
rect 9198 8610 9226 8615
rect 9030 8465 9058 8470
rect 8694 8415 8695 8441
rect 8721 8415 8722 8441
rect 8694 8409 8722 8415
rect 8806 8441 8834 8447
rect 8806 8415 8807 8441
rect 8833 8415 8834 8441
rect 8806 8274 8834 8415
rect 8750 8246 8834 8274
rect 8862 8385 8890 8391
rect 8862 8359 8863 8385
rect 8889 8359 8890 8385
rect 7238 8023 7239 8049
rect 7265 8023 7266 8049
rect 7238 8017 7266 8023
rect 8638 8106 8666 8111
rect 8750 8106 8778 8246
rect 8806 8162 8834 8167
rect 8862 8162 8890 8359
rect 9198 8162 9226 8582
rect 8806 8161 8890 8162
rect 8806 8135 8807 8161
rect 8833 8135 8890 8161
rect 8806 8134 8890 8135
rect 8974 8161 9226 8162
rect 8974 8135 9199 8161
rect 9225 8135 9226 8161
rect 8974 8134 9226 8135
rect 8806 8129 8834 8134
rect 8638 8105 8778 8106
rect 8638 8079 8639 8105
rect 8665 8079 8778 8105
rect 8638 8078 8778 8079
rect 7574 7994 7602 7999
rect 7574 7947 7602 7966
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8638 4214 8666 8078
rect 8974 8049 9002 8134
rect 9198 8129 9226 8134
rect 9254 8442 9282 9870
rect 9310 8666 9338 10038
rect 9422 9897 9450 9903
rect 9422 9871 9423 9897
rect 9449 9871 9450 9897
rect 9366 9842 9394 9847
rect 9366 9673 9394 9814
rect 9366 9647 9367 9673
rect 9393 9647 9394 9673
rect 9366 9641 9394 9647
rect 9422 9170 9450 9871
rect 9478 9898 9506 11159
rect 9590 10906 9618 11550
rect 9534 10289 9562 10295
rect 9534 10263 9535 10289
rect 9561 10263 9562 10289
rect 9534 10066 9562 10263
rect 9590 10094 9618 10878
rect 9702 10458 9730 12502
rect 9870 12474 9898 12479
rect 9870 12417 9898 12446
rect 9870 12391 9871 12417
rect 9897 12391 9898 12417
rect 9870 12385 9898 12391
rect 10094 11858 10122 12727
rect 10150 12642 10178 13455
rect 10486 13258 10514 13263
rect 10598 13258 10626 13263
rect 10486 13257 10598 13258
rect 10486 13231 10487 13257
rect 10513 13231 10598 13257
rect 10486 13230 10598 13231
rect 10486 13225 10514 13230
rect 10598 13225 10626 13230
rect 10430 13145 10458 13151
rect 10430 13119 10431 13145
rect 10457 13119 10458 13145
rect 10150 12609 10178 12614
rect 10206 12753 10234 12759
rect 10206 12727 10207 12753
rect 10233 12727 10234 12753
rect 10206 12698 10234 12727
rect 10374 12754 10402 12759
rect 10374 12707 10402 12726
rect 10206 12586 10234 12670
rect 10206 12553 10234 12558
rect 9814 11830 10122 11858
rect 9758 11242 9786 11247
rect 9758 10962 9786 11214
rect 9814 11186 9842 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10430 11690 10458 13119
rect 10598 13146 10626 13151
rect 10598 12810 10626 13118
rect 10598 12777 10626 12782
rect 10430 11657 10458 11662
rect 10654 12697 10682 13902
rect 10710 13873 10738 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 12446 18746 12474 20600
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 13454 19138 13482 20600
rect 13454 19105 13482 19110
rect 12446 18713 12474 18718
rect 13118 18746 13146 18751
rect 13118 18699 13146 18718
rect 13790 18746 13818 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 14686 19138 14714 19143
rect 14686 19091 14714 19110
rect 13790 18713 13818 18718
rect 14294 19025 14322 19031
rect 14294 18999 14295 19025
rect 14321 18999 14322 19025
rect 12222 15946 12306 15974
rect 12614 18633 12642 18639
rect 12614 18607 12615 18633
rect 12641 18607 12642 18633
rect 12222 14378 12250 15946
rect 12614 15106 12642 18607
rect 14070 18633 14098 18639
rect 14070 18607 14071 18633
rect 14097 18607 14098 18633
rect 14070 15974 14098 18607
rect 12558 15078 12642 15106
rect 13790 15946 14098 15974
rect 12222 14377 12418 14378
rect 12222 14351 12223 14377
rect 12249 14351 12418 14377
rect 12222 14350 12418 14351
rect 12222 14345 12250 14350
rect 10822 14321 10850 14327
rect 10822 14295 10823 14321
rect 10849 14295 10850 14321
rect 10822 14266 10850 14295
rect 10822 14233 10850 14238
rect 11158 14265 11186 14271
rect 11158 14239 11159 14265
rect 11185 14239 11186 14265
rect 11158 14041 11186 14239
rect 11158 14015 11159 14041
rect 11185 14015 11186 14041
rect 11158 14009 11186 14015
rect 12278 14041 12306 14350
rect 12390 14321 12418 14350
rect 12390 14295 12391 14321
rect 12417 14295 12418 14321
rect 12390 14289 12418 14295
rect 12558 14265 12586 15078
rect 12558 14239 12559 14265
rect 12585 14239 12586 14265
rect 12558 14233 12586 14239
rect 12614 14266 12642 14271
rect 12278 14015 12279 14041
rect 12305 14015 12306 14041
rect 12278 14009 12306 14015
rect 11102 13930 11130 13935
rect 11102 13883 11130 13902
rect 11214 13929 11242 13935
rect 11214 13903 11215 13929
rect 11241 13903 11242 13929
rect 10710 13847 10711 13873
rect 10737 13847 10738 13873
rect 10710 13145 10738 13847
rect 10990 13874 11018 13879
rect 10710 13119 10711 13145
rect 10737 13119 10738 13145
rect 10710 13113 10738 13119
rect 10878 13258 10906 13263
rect 10878 12754 10906 13230
rect 10934 12754 10962 12759
rect 10878 12753 10962 12754
rect 10878 12727 10935 12753
rect 10961 12727 10962 12753
rect 10878 12726 10962 12727
rect 10934 12721 10962 12726
rect 10654 12671 10655 12697
rect 10681 12671 10682 12697
rect 9814 11139 9842 11158
rect 9870 11634 9898 11639
rect 9870 11130 9898 11606
rect 10486 11521 10514 11527
rect 10486 11495 10487 11521
rect 10513 11495 10514 11521
rect 9870 11073 9898 11102
rect 9870 11047 9871 11073
rect 9897 11047 9898 11073
rect 9870 11041 9898 11047
rect 10038 11129 10066 11135
rect 10038 11103 10039 11129
rect 10065 11103 10066 11129
rect 10038 11074 10066 11103
rect 10038 11041 10066 11046
rect 10318 11129 10346 11135
rect 10318 11103 10319 11129
rect 10345 11103 10346 11129
rect 10318 11018 10346 11103
rect 10486 11130 10514 11495
rect 10654 11298 10682 12671
rect 10710 12642 10738 12647
rect 10710 12595 10738 12614
rect 10990 12474 11018 13846
rect 11214 13818 11242 13903
rect 11438 13930 11466 13935
rect 11438 13883 11466 13902
rect 12166 13930 12194 13935
rect 12166 13883 12194 13902
rect 12334 13929 12362 13935
rect 12614 13930 12642 14238
rect 12782 14266 12810 14271
rect 12782 14219 12810 14238
rect 12334 13903 12335 13929
rect 12361 13903 12362 13929
rect 12110 13874 12138 13879
rect 11214 13785 11242 13790
rect 12054 13818 12082 13823
rect 12054 13537 12082 13790
rect 12110 13593 12138 13846
rect 12110 13567 12111 13593
rect 12137 13567 12138 13593
rect 12110 13561 12138 13567
rect 12054 13511 12055 13537
rect 12081 13511 12082 13537
rect 12054 13505 12082 13511
rect 11942 13426 11970 13431
rect 11942 13379 11970 13398
rect 12166 13425 12194 13431
rect 12166 13399 12167 13425
rect 12193 13399 12194 13425
rect 11886 13146 11914 13151
rect 11830 12810 11858 12815
rect 11158 12754 11186 12759
rect 11158 12707 11186 12726
rect 11662 12754 11690 12759
rect 11662 12707 11690 12726
rect 10990 12441 11018 12446
rect 11270 12698 11298 12703
rect 11438 12698 11466 12703
rect 11270 12473 11298 12670
rect 11270 12447 11271 12473
rect 11297 12447 11298 12473
rect 11270 12441 11298 12447
rect 11326 12697 11466 12698
rect 11326 12671 11439 12697
rect 11465 12671 11466 12697
rect 11326 12670 11466 12671
rect 10934 12305 10962 12311
rect 10934 12279 10935 12305
rect 10961 12279 10962 12305
rect 10934 12082 10962 12279
rect 10934 12054 11242 12082
rect 11214 12026 11242 12054
rect 11270 12026 11298 12031
rect 11214 12025 11298 12026
rect 11214 11999 11271 12025
rect 11297 11999 11298 12025
rect 11214 11998 11298 11999
rect 11158 11969 11186 11975
rect 11158 11943 11159 11969
rect 11185 11943 11186 11969
rect 10710 11690 10738 11695
rect 10738 11662 10906 11690
rect 10710 11657 10738 11662
rect 10710 11578 10738 11583
rect 10710 11531 10738 11550
rect 10710 11298 10738 11303
rect 10654 11297 10738 11298
rect 10654 11271 10711 11297
rect 10737 11271 10738 11297
rect 10654 11270 10738 11271
rect 10710 11265 10738 11270
rect 10598 11186 10626 11191
rect 10598 11139 10626 11158
rect 10766 11186 10794 11191
rect 10486 11097 10514 11102
rect 9918 10990 10050 10995
rect 10318 10990 10458 11018
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10430 10962 10458 10990
rect 10486 10962 10514 10967
rect 10430 10934 10486 10962
rect 9758 10570 9786 10934
rect 10486 10929 10514 10934
rect 10710 10962 10738 10967
rect 10374 10906 10402 10911
rect 9758 10542 9842 10570
rect 9758 10458 9786 10463
rect 9702 10457 9786 10458
rect 9702 10431 9759 10457
rect 9785 10431 9786 10457
rect 9702 10430 9786 10431
rect 9590 10066 9674 10094
rect 9534 10033 9562 10038
rect 9590 10010 9618 10015
rect 9590 9963 9618 9982
rect 9646 9898 9674 10066
rect 9478 9865 9506 9870
rect 9534 9870 9674 9898
rect 9422 9137 9450 9142
rect 9534 9058 9562 9870
rect 9366 8834 9394 8839
rect 9366 8787 9394 8806
rect 9534 8833 9562 9030
rect 9534 8807 9535 8833
rect 9561 8807 9562 8833
rect 9534 8801 9562 8807
rect 9590 9338 9618 9343
rect 9310 8633 9338 8638
rect 9422 8721 9450 8727
rect 9422 8695 9423 8721
rect 9449 8695 9450 8721
rect 8974 8023 8975 8049
rect 9001 8023 9002 8049
rect 8974 8017 9002 8023
rect 8862 7994 8890 7999
rect 9142 7994 9170 7999
rect 8862 7947 8890 7966
rect 9086 7993 9170 7994
rect 9086 7967 9143 7993
rect 9169 7967 9170 7993
rect 9086 7966 9170 7967
rect 9086 7713 9114 7966
rect 9142 7961 9170 7966
rect 9086 7687 9087 7713
rect 9113 7687 9114 7713
rect 9086 7681 9114 7687
rect 8750 7657 8778 7663
rect 8750 7631 8751 7657
rect 8777 7631 8778 7657
rect 8750 7602 8778 7631
rect 8750 7569 8778 7574
rect 9254 7602 9282 8414
rect 9310 8162 9338 8167
rect 9422 8162 9450 8695
rect 9590 8218 9618 9310
rect 9646 9002 9674 9007
rect 9646 8945 9674 8974
rect 9646 8919 9647 8945
rect 9673 8919 9674 8945
rect 9646 8913 9674 8919
rect 9702 8834 9730 10430
rect 9758 10425 9786 10430
rect 9814 9674 9842 10542
rect 10038 10402 10066 10407
rect 10038 10401 10122 10402
rect 10038 10375 10039 10401
rect 10065 10375 10122 10401
rect 10038 10374 10122 10375
rect 10038 10369 10066 10374
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9814 9627 9842 9646
rect 9870 10122 9898 10127
rect 9870 10065 9898 10094
rect 10094 10122 10122 10374
rect 10094 10089 10122 10094
rect 10150 10401 10178 10407
rect 10150 10375 10151 10401
rect 10177 10375 10178 10401
rect 9870 10039 9871 10065
rect 9897 10039 9898 10065
rect 9870 9617 9898 10039
rect 10150 10010 10178 10375
rect 10150 9977 10178 9982
rect 10206 10122 10234 10127
rect 9926 9842 9954 9847
rect 9926 9674 9954 9814
rect 10094 9786 10122 9791
rect 9926 9641 9954 9646
rect 10038 9730 10066 9735
rect 9870 9591 9871 9617
rect 9897 9591 9898 9617
rect 9870 9585 9898 9591
rect 9758 9561 9786 9567
rect 9758 9535 9759 9561
rect 9785 9535 9786 9561
rect 9758 9338 9786 9535
rect 10038 9562 10066 9702
rect 10094 9673 10122 9758
rect 10206 9730 10234 10094
rect 10374 10065 10402 10878
rect 10430 10402 10458 10407
rect 10654 10402 10682 10407
rect 10430 10401 10682 10402
rect 10430 10375 10431 10401
rect 10457 10375 10655 10401
rect 10681 10375 10682 10401
rect 10430 10374 10682 10375
rect 10430 10290 10458 10374
rect 10654 10369 10682 10374
rect 10430 10257 10458 10262
rect 10710 10094 10738 10934
rect 10374 10039 10375 10065
rect 10401 10039 10402 10065
rect 10374 10033 10402 10039
rect 10654 10066 10738 10094
rect 10766 10122 10794 11158
rect 10878 10094 10906 11662
rect 11046 11634 11074 11639
rect 11046 11633 11130 11634
rect 11046 11607 11047 11633
rect 11073 11607 11130 11633
rect 11046 11606 11130 11607
rect 11046 11601 11074 11606
rect 10934 11242 10962 11247
rect 10934 11195 10962 11214
rect 11046 11242 11074 11247
rect 10094 9647 10095 9673
rect 10121 9647 10122 9673
rect 10094 9641 10122 9647
rect 10150 9702 10234 9730
rect 10038 9529 10066 9534
rect 10094 9562 10122 9567
rect 10150 9562 10178 9702
rect 10374 9617 10402 9623
rect 10374 9591 10375 9617
rect 10401 9591 10402 9617
rect 10094 9561 10178 9562
rect 10094 9535 10095 9561
rect 10121 9535 10178 9561
rect 10094 9534 10178 9535
rect 10206 9562 10234 9567
rect 10094 9529 10122 9534
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10206 9338 10234 9534
rect 9758 9305 9786 9310
rect 10038 9310 10234 9338
rect 9870 9226 9898 9231
rect 9702 8801 9730 8806
rect 9758 8834 9786 8839
rect 9870 8834 9898 9198
rect 10038 9225 10066 9310
rect 10038 9199 10039 9225
rect 10065 9199 10066 9225
rect 10038 9193 10066 9199
rect 10094 9226 10122 9231
rect 10094 9179 10122 9198
rect 10206 9225 10234 9231
rect 10206 9199 10207 9225
rect 10233 9199 10234 9225
rect 10206 9058 10234 9199
rect 10374 9114 10402 9591
rect 10654 9561 10682 10066
rect 10654 9535 10655 9561
rect 10681 9535 10682 9561
rect 10654 9170 10682 9535
rect 10766 9561 10794 10094
rect 10822 10066 10906 10094
rect 10822 9730 10850 10066
rect 10878 9953 10906 9959
rect 10878 9927 10879 9953
rect 10905 9927 10906 9953
rect 10878 9898 10906 9927
rect 10878 9865 10906 9870
rect 10822 9729 10906 9730
rect 10822 9703 10823 9729
rect 10849 9703 10906 9729
rect 10822 9702 10906 9703
rect 10822 9697 10850 9702
rect 10766 9535 10767 9561
rect 10793 9535 10794 9561
rect 10766 9529 10794 9535
rect 10654 9137 10682 9142
rect 10374 9081 10402 9086
rect 10150 8946 10178 8951
rect 10094 8918 10150 8946
rect 10094 8889 10122 8918
rect 10150 8913 10178 8918
rect 10094 8863 10095 8889
rect 10121 8863 10122 8889
rect 10094 8857 10122 8863
rect 10206 8889 10234 9030
rect 10206 8863 10207 8889
rect 10233 8863 10234 8889
rect 10206 8857 10234 8863
rect 10766 9058 10794 9063
rect 9758 8833 9898 8834
rect 9758 8807 9759 8833
rect 9785 8807 9898 8833
rect 9758 8806 9898 8807
rect 10766 8834 10794 9030
rect 9758 8801 9786 8806
rect 10766 8787 10794 8806
rect 10878 8946 10906 9702
rect 11046 9562 11074 11214
rect 11102 10962 11130 11606
rect 11158 11578 11186 11943
rect 11158 11018 11186 11550
rect 11158 10985 11186 10990
rect 11214 11578 11242 11583
rect 11270 11578 11298 11998
rect 11214 11577 11298 11578
rect 11214 11551 11215 11577
rect 11241 11551 11298 11577
rect 11214 11550 11298 11551
rect 11102 10929 11130 10934
rect 11214 10850 11242 11550
rect 11326 11410 11354 12670
rect 11438 12665 11466 12670
rect 11774 12697 11802 12703
rect 11774 12671 11775 12697
rect 11801 12671 11802 12697
rect 11662 12474 11690 12479
rect 11662 12427 11690 12446
rect 11438 12361 11466 12367
rect 11438 12335 11439 12361
rect 11465 12335 11466 12361
rect 11438 12026 11466 12335
rect 11494 12026 11522 12031
rect 11438 12025 11522 12026
rect 11438 11999 11495 12025
rect 11521 11999 11522 12025
rect 11438 11998 11522 11999
rect 11494 11993 11522 11998
rect 11774 11634 11802 12671
rect 11774 11587 11802 11606
rect 11662 11578 11690 11583
rect 11830 11578 11858 12782
rect 11886 12809 11914 13118
rect 11886 12783 11887 12809
rect 11913 12783 11914 12809
rect 11886 12777 11914 12783
rect 11942 13034 11970 13039
rect 11942 12754 11970 13006
rect 12166 12809 12194 13399
rect 12334 13314 12362 13903
rect 12390 13929 12642 13930
rect 12390 13903 12615 13929
rect 12641 13903 12642 13929
rect 12390 13902 12642 13903
rect 12390 13538 12418 13902
rect 12614 13897 12642 13902
rect 13006 13874 13034 13879
rect 13006 13827 13034 13846
rect 12726 13818 12754 13823
rect 12754 13790 12810 13818
rect 12726 13785 12754 13790
rect 12390 13491 12418 13510
rect 12726 13482 12754 13487
rect 12334 13281 12362 13286
rect 12670 13481 12754 13482
rect 12670 13455 12727 13481
rect 12753 13455 12754 13481
rect 12670 13454 12754 13455
rect 12670 13257 12698 13454
rect 12726 13449 12754 13454
rect 12670 13231 12671 13257
rect 12697 13231 12698 13257
rect 12670 13225 12698 13231
rect 12726 13258 12754 13263
rect 12782 13258 12810 13790
rect 13790 13594 13818 15946
rect 14294 14266 14322 18999
rect 14574 18746 14602 18751
rect 14574 18699 14602 18718
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 13510 13593 13818 13594
rect 13510 13567 13791 13593
rect 13817 13567 13818 13593
rect 13510 13566 13818 13567
rect 13174 13538 13202 13543
rect 13118 13426 13146 13431
rect 12726 13257 12810 13258
rect 12726 13231 12727 13257
rect 12753 13231 12810 13257
rect 12726 13230 12810 13231
rect 12894 13314 12922 13319
rect 12726 13225 12754 13230
rect 12614 13146 12642 13151
rect 12614 13099 12642 13118
rect 12166 12783 12167 12809
rect 12193 12783 12194 12809
rect 12166 12777 12194 12783
rect 12054 12754 12082 12759
rect 11942 12753 12082 12754
rect 11942 12727 11943 12753
rect 11969 12727 12055 12753
rect 12081 12727 12082 12753
rect 11942 12726 12082 12727
rect 11942 12721 11970 12726
rect 12054 12721 12082 12726
rect 12222 12753 12250 12759
rect 12222 12727 12223 12753
rect 12249 12727 12250 12753
rect 12166 11634 12194 11639
rect 12222 11634 12250 12727
rect 12390 12698 12418 12703
rect 12390 12651 12418 12670
rect 12894 12473 12922 13286
rect 13118 13257 13146 13398
rect 13118 13231 13119 13257
rect 13145 13231 13146 13257
rect 13118 13225 13146 13231
rect 12950 13146 12978 13151
rect 12950 13099 12978 13118
rect 12894 12447 12895 12473
rect 12921 12447 12922 12473
rect 12894 11970 12922 12447
rect 12894 11937 12922 11942
rect 13062 12361 13090 12367
rect 13062 12335 13063 12361
rect 13089 12335 13090 12361
rect 12194 11606 12250 11634
rect 12670 11858 12698 11863
rect 11886 11578 11914 11583
rect 11662 11577 11746 11578
rect 11662 11551 11663 11577
rect 11689 11551 11746 11577
rect 11662 11550 11746 11551
rect 11830 11577 11914 11578
rect 11830 11551 11887 11577
rect 11913 11551 11914 11577
rect 11830 11550 11914 11551
rect 11662 11545 11690 11550
rect 11326 11382 11466 11410
rect 11382 11242 11410 11247
rect 11382 11195 11410 11214
rect 11214 10817 11242 10822
rect 11326 10794 11354 10799
rect 11326 10747 11354 10766
rect 11214 10010 11242 10015
rect 11214 9963 11242 9982
rect 11438 9730 11466 11382
rect 11662 11242 11690 11247
rect 11718 11242 11746 11550
rect 11886 11545 11914 11550
rect 12054 11577 12082 11583
rect 12054 11551 12055 11577
rect 12081 11551 12082 11577
rect 11998 11466 12026 11471
rect 11942 11465 12026 11466
rect 11942 11439 11999 11465
rect 12025 11439 12026 11465
rect 11942 11438 12026 11439
rect 11774 11242 11802 11247
rect 11718 11241 11802 11242
rect 11718 11215 11775 11241
rect 11801 11215 11802 11241
rect 11718 11214 11802 11215
rect 11494 11130 11522 11135
rect 11494 11083 11522 11102
rect 11662 10905 11690 11214
rect 11662 10879 11663 10905
rect 11689 10879 11690 10905
rect 11662 10873 11690 10879
rect 11774 10906 11802 11214
rect 11550 10850 11578 10855
rect 11774 10850 11802 10878
rect 11830 10850 11858 10855
rect 11774 10849 11858 10850
rect 11774 10823 11831 10849
rect 11857 10823 11858 10849
rect 11774 10822 11858 10823
rect 11550 10793 11578 10822
rect 11830 10817 11858 10822
rect 11550 10767 11551 10793
rect 11577 10767 11578 10793
rect 11550 10761 11578 10767
rect 11774 10738 11802 10743
rect 11046 9529 11074 9534
rect 11326 9729 11466 9730
rect 11326 9703 11439 9729
rect 11465 9703 11466 9729
rect 11326 9702 11466 9703
rect 11214 9225 11242 9231
rect 11214 9199 11215 9225
rect 11241 9199 11242 9225
rect 11102 9169 11130 9175
rect 11102 9143 11103 9169
rect 11129 9143 11130 9169
rect 11046 9114 11074 9119
rect 11046 9067 11074 9086
rect 11102 9002 11130 9143
rect 10878 8833 10906 8918
rect 10990 8974 11130 9002
rect 11158 9114 11186 9119
rect 10990 8945 11018 8974
rect 10990 8919 10991 8945
rect 11017 8919 11018 8945
rect 10990 8913 11018 8919
rect 11102 8890 11130 8895
rect 11158 8890 11186 9086
rect 11214 9058 11242 9199
rect 11214 9025 11242 9030
rect 11102 8889 11186 8890
rect 11102 8863 11103 8889
rect 11129 8863 11186 8889
rect 11102 8862 11186 8863
rect 11102 8857 11130 8862
rect 10878 8807 10879 8833
rect 10905 8807 10906 8833
rect 10878 8801 10906 8807
rect 11214 8778 11242 8783
rect 11214 8777 11298 8778
rect 11214 8751 11215 8777
rect 11241 8751 11298 8777
rect 11214 8750 11298 8751
rect 11214 8745 11242 8750
rect 9926 8722 9954 8741
rect 9926 8689 9954 8694
rect 10934 8721 10962 8727
rect 10934 8695 10935 8721
rect 10961 8695 10962 8721
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10934 8442 10962 8695
rect 11270 8666 11298 8750
rect 11270 8633 11298 8638
rect 10990 8554 11018 8559
rect 10990 8553 11186 8554
rect 10990 8527 10991 8553
rect 11017 8527 11186 8553
rect 10990 8526 11186 8527
rect 10990 8521 11018 8526
rect 11158 8498 11186 8526
rect 11326 8553 11354 9702
rect 11438 9697 11466 9702
rect 11550 10626 11578 10631
rect 11550 9281 11578 10598
rect 11774 10346 11802 10710
rect 11886 10681 11914 10687
rect 11886 10655 11887 10681
rect 11913 10655 11914 10681
rect 11886 10626 11914 10655
rect 11886 10593 11914 10598
rect 11774 10094 11802 10318
rect 11942 10094 11970 11438
rect 11998 11433 12026 11438
rect 11998 11073 12026 11079
rect 11998 11047 11999 11073
rect 12025 11047 12026 11073
rect 11998 11018 12026 11047
rect 12054 11074 12082 11551
rect 12166 11186 12194 11606
rect 12166 11153 12194 11158
rect 12670 11297 12698 11830
rect 12782 11746 12810 11751
rect 12782 11577 12810 11718
rect 13062 11634 13090 12335
rect 13174 12362 13202 13510
rect 13286 13314 13314 13319
rect 13230 13258 13258 13263
rect 13230 13211 13258 13230
rect 13286 13201 13314 13286
rect 13510 13257 13538 13566
rect 13790 13561 13818 13566
rect 14070 14238 14322 14266
rect 14070 13873 14098 14238
rect 14070 13847 14071 13873
rect 14097 13847 14098 13873
rect 14014 13538 14042 13543
rect 14014 13491 14042 13510
rect 13510 13231 13511 13257
rect 13537 13231 13538 13257
rect 13510 13225 13538 13231
rect 13566 13314 13594 13319
rect 13286 13175 13287 13201
rect 13313 13175 13314 13201
rect 13286 13169 13314 13175
rect 13566 13201 13594 13286
rect 14070 13258 14098 13847
rect 14294 13873 14322 13879
rect 14294 13847 14295 13873
rect 14321 13847 14322 13873
rect 14294 13538 14322 13847
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 14294 13505 14322 13510
rect 14910 13538 14938 13543
rect 14070 13225 14098 13230
rect 13566 13175 13567 13201
rect 13593 13175 13594 13201
rect 13566 13169 13594 13175
rect 13398 13146 13426 13151
rect 13398 13099 13426 13118
rect 14910 12473 14938 13510
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 14910 12447 14911 12473
rect 14937 12447 14938 12473
rect 13230 12362 13258 12367
rect 13174 12361 13258 12362
rect 13174 12335 13231 12361
rect 13257 12335 13258 12361
rect 13174 12334 13258 12335
rect 13174 11746 13202 12334
rect 13230 12329 13258 12334
rect 13622 12305 13650 12311
rect 13622 12279 13623 12305
rect 13649 12279 13650 12305
rect 13398 12026 13426 12031
rect 13622 12026 13650 12279
rect 13902 12306 13930 12311
rect 13846 12082 13874 12087
rect 13398 12025 13650 12026
rect 13398 11999 13399 12025
rect 13425 11999 13650 12025
rect 13398 11998 13650 11999
rect 13678 12081 13874 12082
rect 13678 12055 13847 12081
rect 13873 12055 13874 12081
rect 13678 12054 13874 12055
rect 13398 11993 13426 11998
rect 13678 11969 13706 12054
rect 13846 12049 13874 12054
rect 13678 11943 13679 11969
rect 13705 11943 13706 11969
rect 13678 11937 13706 11943
rect 13790 11970 13818 11975
rect 13790 11923 13818 11942
rect 13846 11914 13874 11919
rect 13902 11914 13930 12278
rect 14686 12306 14714 12311
rect 14686 12259 14714 12278
rect 13846 11913 13930 11914
rect 13846 11887 13847 11913
rect 13873 11887 13930 11913
rect 13846 11886 13930 11887
rect 13846 11881 13874 11886
rect 13174 11713 13202 11718
rect 13342 11857 13370 11863
rect 13342 11831 13343 11857
rect 13369 11831 13370 11857
rect 13062 11601 13090 11606
rect 12782 11551 12783 11577
rect 12809 11551 12810 11577
rect 12782 11545 12810 11551
rect 13118 11522 13146 11527
rect 12670 11271 12671 11297
rect 12697 11271 12698 11297
rect 12166 11074 12194 11079
rect 12054 11046 12166 11074
rect 12166 11027 12194 11046
rect 12334 11073 12362 11079
rect 12334 11047 12335 11073
rect 12361 11047 12362 11073
rect 11998 10985 12026 10990
rect 12054 10850 12082 10855
rect 12054 10793 12082 10822
rect 12054 10767 12055 10793
rect 12081 10767 12082 10793
rect 12054 10761 12082 10767
rect 12334 10681 12362 11047
rect 12334 10655 12335 10681
rect 12361 10655 12362 10681
rect 12166 10346 12194 10351
rect 11774 10066 11914 10094
rect 11942 10066 12026 10094
rect 11774 9674 11802 9679
rect 11774 9617 11802 9646
rect 11774 9591 11775 9617
rect 11801 9591 11802 9617
rect 11774 9585 11802 9591
rect 11550 9255 11551 9281
rect 11577 9255 11578 9281
rect 11550 9249 11578 9255
rect 11662 9450 11690 9455
rect 11382 9225 11410 9231
rect 11382 9199 11383 9225
rect 11409 9199 11410 9225
rect 11382 9114 11410 9199
rect 11606 9225 11634 9231
rect 11606 9199 11607 9225
rect 11633 9199 11634 9225
rect 11382 9002 11410 9086
rect 11438 9169 11466 9175
rect 11438 9143 11439 9169
rect 11465 9143 11466 9169
rect 11438 9058 11466 9143
rect 11606 9170 11634 9199
rect 11606 9137 11634 9142
rect 11662 9058 11690 9422
rect 11830 9338 11858 9343
rect 11438 9030 11578 9058
rect 11550 9002 11578 9030
rect 11382 8974 11522 9002
rect 11494 8833 11522 8974
rect 11550 8969 11578 8974
rect 11606 9030 11690 9058
rect 11718 9058 11746 9063
rect 11494 8807 11495 8833
rect 11521 8807 11522 8833
rect 11494 8801 11522 8807
rect 11606 8833 11634 9030
rect 11606 8807 11607 8833
rect 11633 8807 11634 8833
rect 11606 8801 11634 8807
rect 11662 8834 11690 8839
rect 11662 8787 11690 8806
rect 11326 8527 11327 8553
rect 11353 8527 11354 8553
rect 11326 8498 11354 8527
rect 11158 8470 11354 8498
rect 11382 8777 11410 8783
rect 11382 8751 11383 8777
rect 11409 8751 11410 8777
rect 11102 8442 11130 8447
rect 10934 8441 11130 8442
rect 10934 8415 11103 8441
rect 11129 8415 11130 8441
rect 10934 8414 11130 8415
rect 11102 8409 11130 8414
rect 10934 8330 10962 8335
rect 11270 8330 11298 8335
rect 10822 8329 10962 8330
rect 10822 8303 10935 8329
rect 10961 8303 10962 8329
rect 10822 8302 10962 8303
rect 9590 8190 9730 8218
rect 9310 8161 9450 8162
rect 9310 8135 9311 8161
rect 9337 8135 9450 8161
rect 9310 8134 9450 8135
rect 9310 8129 9338 8134
rect 9646 8106 9674 8111
rect 9422 8105 9674 8106
rect 9422 8079 9647 8105
rect 9673 8079 9674 8105
rect 9422 8078 9674 8079
rect 9422 8049 9450 8078
rect 9646 8073 9674 8078
rect 9422 8023 9423 8049
rect 9449 8023 9450 8049
rect 9422 8017 9450 8023
rect 9590 7994 9618 7999
rect 9702 7994 9730 8190
rect 9590 7993 9730 7994
rect 9590 7967 9591 7993
rect 9617 7967 9730 7993
rect 9590 7966 9730 7967
rect 9758 8049 9786 8055
rect 9758 8023 9759 8049
rect 9785 8023 9786 8049
rect 9590 7961 9618 7966
rect 9254 7569 9282 7574
rect 9758 7490 9786 8023
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 10822 7713 10850 8302
rect 10934 8297 10962 8302
rect 11158 8329 11298 8330
rect 11158 8303 11271 8329
rect 11297 8303 11298 8329
rect 11158 8302 11298 8303
rect 10822 7687 10823 7713
rect 10849 7687 10850 7713
rect 10822 7681 10850 7687
rect 10486 7657 10514 7663
rect 10486 7631 10487 7657
rect 10513 7631 10514 7657
rect 10150 7602 10178 7607
rect 9982 7601 10178 7602
rect 9982 7575 10151 7601
rect 10177 7575 10178 7601
rect 9982 7574 10178 7575
rect 9982 7490 10010 7574
rect 10150 7569 10178 7574
rect 10318 7602 10346 7607
rect 9758 7462 10010 7490
rect 8638 4186 8834 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8750 1834 8778 1839
rect 8750 400 8778 1806
rect 8806 1777 8834 4186
rect 9814 2170 9842 7462
rect 10318 7321 10346 7574
rect 10486 7602 10514 7631
rect 10486 7569 10514 7574
rect 10318 7295 10319 7321
rect 10345 7295 10346 7321
rect 10318 7289 10346 7295
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 11158 6929 11186 8302
rect 11270 8297 11298 8302
rect 11158 6903 11159 6929
rect 11185 6903 11186 6929
rect 11158 6897 11186 6903
rect 10094 6818 10122 6823
rect 10094 6771 10122 6790
rect 10710 6818 10738 6823
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9870 2170 9898 2175
rect 9814 2169 9898 2170
rect 9814 2143 9871 2169
rect 9897 2143 9898 2169
rect 9814 2142 9898 2143
rect 9870 2137 9898 2142
rect 9758 2058 9786 2063
rect 9310 1834 9338 1839
rect 9310 1787 9338 1806
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9758 400 9786 2030
rect 10374 2058 10402 2063
rect 10374 2011 10402 2030
rect 10710 1777 10738 6790
rect 11382 6818 11410 8751
rect 11550 8721 11578 8727
rect 11550 8695 11551 8721
rect 11577 8695 11578 8721
rect 11550 8554 11578 8695
rect 11438 8526 11578 8554
rect 11606 8666 11634 8671
rect 11438 8497 11466 8526
rect 11438 8471 11439 8497
rect 11465 8471 11466 8497
rect 11438 8465 11466 8471
rect 11606 7602 11634 8638
rect 11662 8554 11690 8559
rect 11718 8554 11746 9030
rect 11662 8553 11746 8554
rect 11662 8527 11663 8553
rect 11689 8527 11746 8553
rect 11662 8526 11746 8527
rect 11662 8521 11690 8526
rect 11830 8498 11858 9310
rect 11886 8777 11914 10066
rect 11998 9225 12026 10066
rect 12054 10009 12082 10015
rect 12054 9983 12055 10009
rect 12081 9983 12082 10009
rect 12054 9674 12082 9983
rect 12054 9641 12082 9646
rect 12110 9898 12138 9903
rect 12110 9617 12138 9870
rect 12110 9591 12111 9617
rect 12137 9591 12138 9617
rect 12110 9562 12138 9591
rect 12110 9529 12138 9534
rect 12166 9394 12194 10318
rect 12222 10066 12250 10071
rect 12222 10019 12250 10038
rect 12334 10010 12362 10655
rect 12614 10794 12642 10799
rect 12614 10457 12642 10766
rect 12614 10431 12615 10457
rect 12641 10431 12642 10457
rect 12614 10425 12642 10431
rect 12670 10066 12698 11271
rect 13006 11521 13146 11522
rect 13006 11495 13119 11521
rect 13145 11495 13146 11521
rect 13006 11494 13146 11495
rect 13006 11297 13034 11494
rect 13118 11489 13146 11494
rect 13006 11271 13007 11297
rect 13033 11271 13034 11297
rect 13006 11265 13034 11271
rect 12782 11186 12810 11191
rect 12670 10033 12698 10038
rect 12726 11185 12810 11186
rect 12726 11159 12783 11185
rect 12809 11159 12810 11185
rect 12726 11158 12810 11159
rect 12726 11074 12754 11158
rect 12782 11153 12810 11158
rect 12950 11186 12978 11191
rect 12950 11139 12978 11158
rect 13286 11185 13314 11191
rect 13286 11159 13287 11185
rect 13313 11159 13314 11185
rect 13062 11130 13090 11135
rect 13062 11083 13090 11102
rect 12222 9618 12250 9623
rect 12222 9571 12250 9590
rect 12334 9617 12362 9982
rect 12334 9591 12335 9617
rect 12361 9591 12362 9617
rect 12334 9585 12362 9591
rect 11998 9199 11999 9225
rect 12025 9199 12026 9225
rect 11998 9193 12026 9199
rect 12054 9366 12194 9394
rect 12502 9562 12530 9567
rect 12054 9114 12082 9366
rect 12222 9225 12250 9231
rect 12222 9199 12223 9225
rect 12249 9199 12250 9225
rect 12110 9170 12138 9175
rect 12110 9123 12138 9142
rect 11942 9002 11970 9007
rect 11970 8974 12026 9002
rect 11942 8969 11970 8974
rect 11886 8751 11887 8777
rect 11913 8751 11914 8777
rect 11886 8745 11914 8751
rect 11998 8554 12026 8974
rect 12054 8833 12082 9086
rect 12054 8807 12055 8833
rect 12081 8807 12082 8833
rect 12054 8801 12082 8807
rect 12054 8554 12082 8559
rect 11998 8553 12082 8554
rect 11998 8527 12055 8553
rect 12081 8527 12082 8553
rect 11998 8526 12082 8527
rect 12054 8521 12082 8526
rect 11942 8498 11970 8503
rect 11830 8497 11970 8498
rect 11830 8471 11943 8497
rect 11969 8471 11970 8497
rect 11830 8470 11970 8471
rect 11942 8465 11970 8470
rect 12166 8498 12194 8503
rect 12166 8451 12194 8470
rect 11718 8386 11746 8391
rect 11718 8339 11746 8358
rect 12110 8385 12138 8391
rect 12110 8359 12111 8385
rect 12137 8359 12138 8385
rect 11774 8330 11802 8335
rect 12110 8330 12138 8359
rect 11774 8329 12138 8330
rect 11774 8303 11775 8329
rect 11801 8303 12138 8329
rect 11774 8302 12138 8303
rect 11774 8297 11802 8302
rect 12222 8162 12250 9199
rect 12334 9225 12362 9231
rect 12334 9199 12335 9225
rect 12361 9199 12362 9225
rect 12278 9114 12306 9119
rect 12278 8441 12306 9086
rect 12334 9058 12362 9199
rect 12362 9030 12418 9058
rect 12334 9025 12362 9030
rect 12390 8833 12418 9030
rect 12390 8807 12391 8833
rect 12417 8807 12418 8833
rect 12390 8801 12418 8807
rect 12502 8833 12530 9534
rect 12726 9450 12754 11046
rect 12838 11018 12866 11023
rect 12838 10178 12866 10990
rect 12838 9953 12866 10150
rect 13286 10094 13314 11159
rect 13342 10738 13370 11831
rect 13454 11858 13482 11863
rect 13454 11811 13482 11830
rect 14406 11690 14434 11695
rect 13734 11634 13762 11639
rect 13398 11242 13426 11247
rect 13398 11195 13426 11214
rect 13622 11185 13650 11191
rect 13622 11159 13623 11185
rect 13649 11159 13650 11185
rect 13510 11130 13538 11135
rect 13342 10705 13370 10710
rect 13454 11129 13538 11130
rect 13454 11103 13511 11129
rect 13537 11103 13538 11129
rect 13454 11102 13538 11103
rect 13398 10346 13426 10351
rect 13398 10299 13426 10318
rect 13454 10094 13482 11102
rect 13510 11097 13538 11102
rect 13622 10626 13650 11159
rect 13622 10593 13650 10598
rect 13678 11129 13706 11135
rect 13678 11103 13679 11129
rect 13705 11103 13706 11129
rect 13678 10401 13706 11103
rect 13678 10375 13679 10401
rect 13705 10375 13706 10401
rect 13678 10369 13706 10375
rect 13734 11130 13762 11606
rect 13902 11578 13930 11583
rect 13846 11130 13874 11135
rect 13734 11129 13874 11130
rect 13734 11103 13847 11129
rect 13873 11103 13874 11129
rect 13734 11102 13874 11103
rect 13734 10402 13762 11102
rect 13846 11097 13874 11102
rect 13902 11129 13930 11550
rect 14182 11578 14210 11583
rect 14182 11521 14210 11550
rect 14182 11495 14183 11521
rect 14209 11495 14210 11521
rect 14182 11489 14210 11495
rect 13902 11103 13903 11129
rect 13929 11103 13930 11129
rect 13902 11097 13930 11103
rect 14014 11130 14042 11135
rect 14014 11083 14042 11102
rect 14406 10850 14434 11662
rect 14910 11690 14938 12447
rect 18830 12753 18858 12759
rect 18830 12727 18831 12753
rect 18857 12727 18858 12753
rect 18830 12306 18858 12727
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 18830 12273 18858 12278
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 14910 11657 14938 11662
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 14406 10849 14546 10850
rect 14406 10823 14407 10849
rect 14433 10823 14546 10849
rect 14406 10822 14546 10823
rect 14406 10817 14434 10822
rect 13734 10369 13762 10374
rect 13790 10794 13818 10799
rect 14294 10794 14322 10799
rect 13566 10346 13594 10351
rect 13566 10299 13594 10318
rect 13790 10345 13818 10766
rect 14238 10766 14294 10794
rect 13902 10626 13930 10631
rect 13846 10402 13874 10407
rect 13846 10355 13874 10374
rect 13790 10319 13791 10345
rect 13817 10319 13818 10345
rect 13790 10313 13818 10319
rect 13510 10290 13538 10295
rect 13510 10243 13538 10262
rect 13286 10066 13370 10094
rect 13286 10033 13314 10038
rect 12838 9927 12839 9953
rect 12865 9927 12866 9953
rect 12838 9921 12866 9927
rect 13230 9618 13258 9623
rect 13230 9571 13258 9590
rect 13342 9618 13370 10066
rect 13342 9585 13370 9590
rect 13398 10066 13482 10094
rect 13286 9506 13314 9511
rect 12726 9417 12754 9422
rect 13118 9505 13314 9506
rect 13118 9479 13287 9505
rect 13313 9479 13314 9505
rect 13118 9478 13314 9479
rect 12614 9226 12642 9231
rect 12614 9179 12642 9198
rect 12838 9225 12866 9231
rect 12838 9199 12839 9225
rect 12865 9199 12866 9225
rect 12670 9114 12698 9119
rect 12670 9067 12698 9086
rect 12502 8807 12503 8833
rect 12529 8807 12530 8833
rect 12502 8801 12530 8807
rect 12726 8833 12754 8839
rect 12838 8834 12866 9199
rect 13118 9058 13146 9478
rect 13286 9473 13314 9478
rect 13342 9505 13370 9511
rect 13342 9479 13343 9505
rect 13369 9479 13370 9505
rect 13342 9450 13370 9479
rect 13342 9417 13370 9422
rect 13230 9226 13258 9231
rect 13398 9226 13426 10066
rect 13902 10065 13930 10598
rect 13902 10039 13903 10065
rect 13929 10039 13930 10065
rect 13902 10033 13930 10039
rect 14238 9898 14266 10766
rect 14294 10761 14322 10766
rect 14518 10122 14546 10822
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10681 20034 10687
rect 20006 10655 20007 10681
rect 20033 10655 20034 10681
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10458 20034 10655
rect 20006 10425 20034 10430
rect 14294 10121 14546 10122
rect 14294 10095 14519 10121
rect 14545 10095 14546 10121
rect 14294 10094 14546 10095
rect 14294 10009 14322 10094
rect 14294 9983 14295 10009
rect 14321 9983 14322 10009
rect 14294 9977 14322 9983
rect 14238 9870 14322 9898
rect 13510 9618 13538 9623
rect 13510 9571 13538 9590
rect 13230 9225 13426 9226
rect 13230 9199 13231 9225
rect 13257 9199 13426 9225
rect 13230 9198 13426 9199
rect 13230 9193 13258 9198
rect 13118 9025 13146 9030
rect 13174 9170 13202 9175
rect 12726 8807 12727 8833
rect 12753 8807 12754 8833
rect 12614 8778 12642 8783
rect 12614 8731 12642 8750
rect 12278 8415 12279 8441
rect 12305 8415 12306 8441
rect 12278 8409 12306 8415
rect 12222 8129 12250 8134
rect 12558 8386 12586 8391
rect 12558 8105 12586 8358
rect 12558 8079 12559 8105
rect 12585 8079 12586 8105
rect 12558 8073 12586 8079
rect 12166 8050 12194 8055
rect 11998 8022 12166 8050
rect 11662 7602 11690 7607
rect 11606 7574 11662 7602
rect 11662 7569 11690 7574
rect 11886 7602 11914 7607
rect 11886 7555 11914 7574
rect 11494 7546 11522 7551
rect 11494 6930 11522 7518
rect 11998 7153 12026 8022
rect 12166 8003 12194 8022
rect 12726 7938 12754 8807
rect 12782 8833 12866 8834
rect 12782 8807 12839 8833
rect 12865 8807 12866 8833
rect 12782 8806 12866 8807
rect 12782 8442 12810 8806
rect 12838 8801 12866 8806
rect 13174 8497 13202 9142
rect 14294 9169 14322 9870
rect 14518 9338 14546 10094
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 14518 9337 14658 9338
rect 14518 9311 14519 9337
rect 14545 9311 14658 9337
rect 14518 9310 14658 9311
rect 14518 9305 14546 9310
rect 14294 9143 14295 9169
rect 14321 9143 14322 9169
rect 14294 9137 14322 9143
rect 13398 9114 13426 9119
rect 13342 8890 13370 8895
rect 13230 8778 13258 8783
rect 13230 8731 13258 8750
rect 13174 8471 13175 8497
rect 13201 8471 13202 8497
rect 13174 8465 13202 8471
rect 12782 8050 12810 8414
rect 12782 8017 12810 8022
rect 12726 7910 13258 7938
rect 13230 7769 13258 7910
rect 13230 7743 13231 7769
rect 13257 7743 13258 7769
rect 13230 7737 13258 7743
rect 13342 7769 13370 8862
rect 13342 7743 13343 7769
rect 13369 7743 13370 7769
rect 13342 7737 13370 7743
rect 13398 8050 13426 9086
rect 14294 8890 14322 8895
rect 14630 8890 14658 9310
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 14294 8722 14322 8862
rect 14294 8689 14322 8694
rect 14462 8889 14658 8890
rect 14462 8863 14631 8889
rect 14657 8863 14658 8889
rect 14462 8862 14658 8863
rect 14462 8554 14490 8862
rect 14630 8857 14658 8862
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 18886 8833 18914 8839
rect 18886 8807 18887 8833
rect 18913 8807 18914 8833
rect 14126 8553 14490 8554
rect 14126 8527 14463 8553
rect 14489 8527 14490 8553
rect 14126 8526 14490 8527
rect 13622 8498 13650 8503
rect 13622 8106 13650 8470
rect 14126 8442 14154 8526
rect 14462 8521 14490 8526
rect 18830 8722 18858 8727
rect 13958 8386 13986 8391
rect 13902 8358 13958 8386
rect 13846 8162 13874 8167
rect 13846 8115 13874 8134
rect 13622 8059 13650 8078
rect 11998 7127 11999 7153
rect 12025 7127 12026 7153
rect 11494 6873 11522 6902
rect 11774 6930 11802 6935
rect 11998 6930 12026 7127
rect 11802 6902 12026 6930
rect 12054 7713 12082 7719
rect 12054 7687 12055 7713
rect 12081 7687 12082 7713
rect 11774 6883 11802 6902
rect 11494 6847 11495 6873
rect 11521 6847 11522 6873
rect 11494 6841 11522 6847
rect 11382 6785 11410 6790
rect 12054 4214 12082 7687
rect 13398 7713 13426 8022
rect 13790 8050 13818 8055
rect 13790 8003 13818 8022
rect 13846 7994 13874 7999
rect 13902 7994 13930 8358
rect 13958 8353 13986 8358
rect 14126 8105 14154 8414
rect 18830 8441 18858 8694
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 18830 8409 18858 8415
rect 14238 8386 14266 8391
rect 14238 8339 14266 8358
rect 18886 8386 18914 8807
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 18886 8353 18914 8358
rect 20006 8442 20034 8447
rect 20006 8385 20034 8414
rect 20006 8359 20007 8385
rect 20033 8359 20034 8385
rect 20006 8353 20034 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 14126 8079 14127 8105
rect 14153 8079 14154 8105
rect 14126 8073 14154 8079
rect 18830 8106 18858 8111
rect 18830 8049 18858 8078
rect 20006 8106 20034 8111
rect 20006 8059 20034 8078
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 18830 8017 18858 8023
rect 13846 7993 13930 7994
rect 13846 7967 13847 7993
rect 13873 7967 13930 7993
rect 13846 7966 13930 7967
rect 13846 7961 13874 7966
rect 13398 7687 13399 7713
rect 13425 7687 13426 7713
rect 13398 7681 13426 7687
rect 11886 4186 12082 4214
rect 12222 7657 12250 7663
rect 12222 7631 12223 7657
rect 12249 7631 12250 7657
rect 12222 7602 12250 7631
rect 12222 4214 12250 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 12222 4186 12306 4214
rect 11774 2618 11802 2623
rect 10710 1751 10711 1777
rect 10737 1751 10738 1777
rect 10710 1745 10738 1751
rect 11438 1834 11466 1839
rect 11214 1666 11242 1671
rect 11102 1665 11242 1666
rect 11102 1639 11215 1665
rect 11241 1639 11242 1665
rect 11102 1638 11242 1639
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 11102 400 11130 1638
rect 11214 1633 11242 1638
rect 11438 400 11466 1806
rect 11774 400 11802 2590
rect 11886 2561 11914 4186
rect 11886 2535 11887 2561
rect 11913 2535 11914 2561
rect 11886 2529 11914 2535
rect 12278 1777 12306 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12390 2618 12418 2623
rect 12390 2571 12418 2590
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 8736 0 8792 400
rect 9744 0 9800 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 10766 19110 10794 19138
rect 11214 19137 11242 19138
rect 11214 19111 11215 19137
rect 11215 19111 11241 19137
rect 11241 19111 11242 19137
rect 11214 19110 11242 19111
rect 12110 19110 12138 19138
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 854 18185 882 18186
rect 854 18159 855 18185
rect 855 18159 881 18185
rect 881 18159 882 18185
rect 854 18158 882 18159
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2086 14126 2114 14154
rect 966 13454 994 13482
rect 1022 13118 1050 13146
rect 966 12782 994 12810
rect 966 11774 994 11802
rect 966 10430 994 10458
rect 2142 13929 2170 13930
rect 2142 13903 2143 13929
rect 2143 13903 2169 13929
rect 2169 13903 2170 13929
rect 2142 13902 2170 13903
rect 7630 13902 7658 13930
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2142 13537 2170 13538
rect 2142 13511 2143 13537
rect 2143 13511 2169 13537
rect 2169 13511 2170 13537
rect 2142 13510 2170 13511
rect 7294 13510 7322 13538
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 5950 13118 5978 13146
rect 8918 13790 8946 13818
rect 7462 13118 7490 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 7406 13062 7434 13090
rect 6958 12446 6986 12474
rect 7742 13145 7770 13146
rect 7742 13119 7743 13145
rect 7743 13119 7769 13145
rect 7769 13119 7770 13145
rect 7742 13118 7770 13119
rect 8694 13145 8722 13146
rect 8694 13119 8695 13145
rect 8695 13119 8721 13145
rect 8721 13119 8722 13145
rect 8694 13118 8722 13119
rect 7630 13062 7658 13090
rect 8022 13089 8050 13090
rect 8022 13063 8023 13089
rect 8023 13063 8049 13089
rect 8049 13063 8050 13089
rect 8022 13062 8050 13063
rect 7966 12809 7994 12810
rect 7966 12783 7967 12809
rect 7967 12783 7993 12809
rect 7993 12783 7994 12809
rect 7966 12782 7994 12783
rect 8750 12782 8778 12810
rect 7798 12502 7826 12530
rect 7742 12473 7770 12474
rect 7742 12447 7743 12473
rect 7743 12447 7769 12473
rect 7769 12447 7770 12473
rect 7742 12446 7770 12447
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 10654 13902 10682 13930
rect 9366 13846 9394 13874
rect 8806 12502 8834 12530
rect 7910 12446 7938 12474
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 5558 11942 5586 11970
rect 6846 11942 6874 11970
rect 6902 11913 6930 11914
rect 6902 11887 6903 11913
rect 6903 11887 6929 11913
rect 6929 11887 6930 11913
rect 6902 11886 6930 11887
rect 6622 11689 6650 11690
rect 6622 11663 6623 11689
rect 6623 11663 6649 11689
rect 6649 11663 6650 11689
rect 6622 11662 6650 11663
rect 9142 13118 9170 13146
rect 9030 13006 9058 13034
rect 9198 13006 9226 13034
rect 9310 13006 9338 13034
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9366 13062 9394 13090
rect 9534 13006 9562 13034
rect 9086 12446 9114 12474
rect 7742 11913 7770 11914
rect 7742 11887 7743 11913
rect 7743 11887 7769 11913
rect 7769 11887 7770 11913
rect 7742 11886 7770 11887
rect 7238 11830 7266 11858
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6566 10905 6594 10906
rect 6566 10879 6567 10905
rect 6567 10879 6593 10905
rect 6593 10879 6594 10905
rect 6566 10878 6594 10879
rect 2142 10793 2170 10794
rect 2142 10767 2143 10793
rect 2143 10767 2169 10793
rect 2169 10767 2170 10793
rect 2142 10766 2170 10767
rect 4998 10766 5026 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 4998 10457 5026 10458
rect 4998 10431 4999 10457
rect 4999 10431 5025 10457
rect 5025 10431 5026 10457
rect 4998 10430 5026 10431
rect 6678 10430 6706 10458
rect 2086 10262 2114 10290
rect 6398 10065 6426 10066
rect 6398 10039 6399 10065
rect 6399 10039 6425 10065
rect 6425 10039 6426 10065
rect 6398 10038 6426 10039
rect 6902 10878 6930 10906
rect 8022 11857 8050 11858
rect 8022 11831 8023 11857
rect 8023 11831 8049 11857
rect 8049 11831 8050 11857
rect 8022 11830 8050 11831
rect 8078 11662 8106 11690
rect 8190 11662 8218 11690
rect 8302 11158 8330 11186
rect 8414 10905 8442 10906
rect 8414 10879 8415 10905
rect 8415 10879 8441 10905
rect 8441 10879 8442 10905
rect 8414 10878 8442 10879
rect 8470 10822 8498 10850
rect 8302 10793 8330 10794
rect 8302 10767 8303 10793
rect 8303 10767 8329 10793
rect 8329 10767 8330 10793
rect 8302 10766 8330 10767
rect 7910 10486 7938 10514
rect 7966 10374 7994 10402
rect 7798 10206 7826 10234
rect 7742 10094 7770 10122
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6734 9254 6762 9282
rect 2142 9225 2170 9226
rect 2142 9199 2143 9225
rect 2143 9199 2169 9225
rect 2169 9199 2170 9225
rect 2142 9198 2170 9199
rect 5446 9198 5474 9226
rect 7182 10065 7210 10066
rect 7182 10039 7183 10065
rect 7183 10039 7209 10065
rect 7209 10039 7210 10065
rect 7182 10038 7210 10039
rect 7238 10009 7266 10010
rect 7238 9983 7239 10009
rect 7239 9983 7265 10009
rect 7265 9983 7266 10009
rect 7238 9982 7266 9983
rect 7574 10009 7602 10010
rect 7574 9983 7575 10009
rect 7575 9983 7601 10009
rect 7601 9983 7602 10009
rect 7574 9982 7602 9983
rect 7910 10009 7938 10010
rect 7910 9983 7911 10009
rect 7911 9983 7937 10009
rect 7937 9983 7938 10009
rect 7910 9982 7938 9983
rect 7182 9758 7210 9786
rect 966 9113 994 9114
rect 966 9087 967 9113
rect 967 9087 993 9113
rect 993 9087 994 9113
rect 966 9086 994 9087
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 6342 8806 6370 8834
rect 966 8414 994 8442
rect 6902 9142 6930 9170
rect 7182 9281 7210 9282
rect 7182 9255 7183 9281
rect 7183 9255 7209 9281
rect 7209 9255 7210 9281
rect 7182 9254 7210 9255
rect 7126 9198 7154 9226
rect 7406 9169 7434 9170
rect 7406 9143 7407 9169
rect 7407 9143 7433 9169
rect 7433 9143 7434 9169
rect 7406 9142 7434 9143
rect 7238 8777 7266 8778
rect 7238 8751 7239 8777
rect 7239 8751 7265 8777
rect 7265 8751 7266 8777
rect 7238 8750 7266 8751
rect 6846 8694 6874 8722
rect 7238 8414 7266 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 8078 10065 8106 10066
rect 8078 10039 8079 10065
rect 8079 10039 8105 10065
rect 8105 10039 8106 10065
rect 8078 10038 8106 10039
rect 8638 11689 8666 11690
rect 8638 11663 8639 11689
rect 8639 11663 8665 11689
rect 8665 11663 8666 11689
rect 8638 11662 8666 11663
rect 8750 11689 8778 11690
rect 8750 11663 8751 11689
rect 8751 11663 8777 11689
rect 8777 11663 8778 11689
rect 8750 11662 8778 11663
rect 8582 10513 8610 10514
rect 8582 10487 8583 10513
rect 8583 10487 8609 10513
rect 8609 10487 8610 10513
rect 8582 10486 8610 10487
rect 8582 10401 8610 10402
rect 8582 10375 8583 10401
rect 8583 10375 8609 10401
rect 8609 10375 8610 10401
rect 8582 10374 8610 10375
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9646 12502 9674 12530
rect 9310 11689 9338 11690
rect 9310 11663 9311 11689
rect 9311 11663 9337 11689
rect 9337 11663 9338 11689
rect 9310 11662 9338 11663
rect 8694 10206 8722 10234
rect 9086 11185 9114 11186
rect 9086 11159 9087 11185
rect 9087 11159 9113 11185
rect 9113 11159 9114 11185
rect 9086 11158 9114 11159
rect 9310 11158 9338 11186
rect 9422 10934 9450 10962
rect 8806 10849 8834 10850
rect 8806 10823 8807 10849
rect 8807 10823 8833 10849
rect 8833 10823 8834 10849
rect 8806 10822 8834 10823
rect 9142 10822 9170 10850
rect 8750 10766 8778 10794
rect 8246 10094 8274 10122
rect 8750 10094 8778 10122
rect 9086 10374 9114 10402
rect 8190 9982 8218 10010
rect 8246 9926 8274 9954
rect 8134 8806 8162 8834
rect 8078 8777 8106 8778
rect 8078 8751 8079 8777
rect 8079 8751 8105 8777
rect 8105 8751 8106 8777
rect 8078 8750 8106 8751
rect 8246 8833 8274 8834
rect 8246 8807 8247 8833
rect 8247 8807 8273 8833
rect 8273 8807 8274 8833
rect 8246 8806 8274 8807
rect 8862 10038 8890 10066
rect 8806 10009 8834 10010
rect 8806 9983 8807 10009
rect 8807 9983 8833 10009
rect 8833 9983 8834 10009
rect 8806 9982 8834 9983
rect 8974 10009 9002 10010
rect 8974 9983 8975 10009
rect 8975 9983 9001 10009
rect 9001 9983 9002 10009
rect 8974 9982 9002 9983
rect 8414 9310 8442 9338
rect 8414 9225 8442 9226
rect 8414 9199 8415 9225
rect 8415 9199 8441 9225
rect 8441 9199 8442 9225
rect 8414 9198 8442 9199
rect 8750 9198 8778 9226
rect 8918 9310 8946 9338
rect 8974 9225 9002 9226
rect 8974 9199 8975 9225
rect 8975 9199 9001 9225
rect 9001 9199 9002 9225
rect 8974 9198 9002 9199
rect 9142 10065 9170 10066
rect 9142 10039 9143 10065
rect 9143 10039 9169 10065
rect 9169 10039 9170 10065
rect 9142 10038 9170 10039
rect 9142 9870 9170 9898
rect 9310 10318 9338 10346
rect 9310 10206 9338 10234
rect 9254 10094 9282 10122
rect 9198 9534 9226 9562
rect 8302 8777 8330 8778
rect 8302 8751 8303 8777
rect 8303 8751 8329 8777
rect 8329 8751 8330 8777
rect 8302 8750 8330 8751
rect 8694 8750 8722 8778
rect 7462 8414 7490 8442
rect 7798 8441 7826 8442
rect 7798 8415 7799 8441
rect 7799 8415 7825 8441
rect 7825 8415 7826 8441
rect 7798 8414 7826 8415
rect 8022 8441 8050 8442
rect 8022 8415 8023 8441
rect 8023 8415 8049 8441
rect 8049 8415 8050 8441
rect 8022 8414 8050 8415
rect 9142 9086 9170 9114
rect 8918 8721 8946 8722
rect 8918 8695 8919 8721
rect 8919 8695 8945 8721
rect 8945 8695 8946 8721
rect 8918 8694 8946 8695
rect 9198 8806 9226 8834
rect 9142 8750 9170 8778
rect 9198 8694 9226 8722
rect 9198 8582 9226 8610
rect 7574 7993 7602 7994
rect 7574 7967 7575 7993
rect 7575 7967 7601 7993
rect 7601 7967 7602 7993
rect 7574 7966 7602 7967
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 9366 9814 9394 9842
rect 9590 10878 9618 10906
rect 9870 12446 9898 12474
rect 10598 13230 10626 13258
rect 10150 12614 10178 12642
rect 10374 12753 10402 12754
rect 10374 12727 10375 12753
rect 10375 12727 10401 12753
rect 10401 12727 10402 12753
rect 10374 12726 10402 12727
rect 10206 12670 10234 12698
rect 10206 12558 10234 12586
rect 9758 11214 9786 11242
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10598 13145 10626 13146
rect 10598 13119 10599 13145
rect 10599 13119 10625 13145
rect 10625 13119 10626 13145
rect 10598 13118 10626 13119
rect 10598 12782 10626 12810
rect 10430 11662 10458 11690
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 13454 19110 13482 19138
rect 12446 18718 12474 18746
rect 13118 18745 13146 18746
rect 13118 18719 13119 18745
rect 13119 18719 13145 18745
rect 13145 18719 13146 18745
rect 13118 18718 13146 18719
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 14686 19137 14714 19138
rect 14686 19111 14687 19137
rect 14687 19111 14713 19137
rect 14713 19111 14714 19137
rect 14686 19110 14714 19111
rect 13790 18718 13818 18746
rect 10822 14238 10850 14266
rect 12614 14238 12642 14266
rect 11102 13929 11130 13930
rect 11102 13903 11103 13929
rect 11103 13903 11129 13929
rect 11129 13903 11130 13929
rect 11102 13902 11130 13903
rect 10990 13873 11018 13874
rect 10990 13847 10991 13873
rect 10991 13847 11017 13873
rect 11017 13847 11018 13873
rect 10990 13846 11018 13847
rect 10878 13230 10906 13258
rect 9814 11185 9842 11186
rect 9814 11159 9815 11185
rect 9815 11159 9841 11185
rect 9841 11159 9842 11185
rect 9814 11158 9842 11159
rect 9870 11606 9898 11634
rect 9870 11102 9898 11130
rect 10038 11046 10066 11074
rect 10710 12641 10738 12642
rect 10710 12615 10711 12641
rect 10711 12615 10737 12641
rect 10737 12615 10738 12641
rect 10710 12614 10738 12615
rect 11438 13929 11466 13930
rect 11438 13903 11439 13929
rect 11439 13903 11465 13929
rect 11465 13903 11466 13929
rect 11438 13902 11466 13903
rect 12166 13929 12194 13930
rect 12166 13903 12167 13929
rect 12167 13903 12193 13929
rect 12193 13903 12194 13929
rect 12166 13902 12194 13903
rect 12782 14265 12810 14266
rect 12782 14239 12783 14265
rect 12783 14239 12809 14265
rect 12809 14239 12810 14265
rect 12782 14238 12810 14239
rect 12110 13846 12138 13874
rect 11214 13790 11242 13818
rect 12054 13790 12082 13818
rect 11942 13425 11970 13426
rect 11942 13399 11943 13425
rect 11943 13399 11969 13425
rect 11969 13399 11970 13425
rect 11942 13398 11970 13399
rect 11886 13118 11914 13146
rect 11830 12782 11858 12810
rect 11158 12753 11186 12754
rect 11158 12727 11159 12753
rect 11159 12727 11185 12753
rect 11185 12727 11186 12753
rect 11158 12726 11186 12727
rect 11662 12753 11690 12754
rect 11662 12727 11663 12753
rect 11663 12727 11689 12753
rect 11689 12727 11690 12753
rect 11662 12726 11690 12727
rect 10990 12446 11018 12474
rect 11270 12670 11298 12698
rect 10710 11662 10738 11690
rect 10710 11577 10738 11578
rect 10710 11551 10711 11577
rect 10711 11551 10737 11577
rect 10737 11551 10738 11577
rect 10710 11550 10738 11551
rect 10598 11185 10626 11186
rect 10598 11159 10599 11185
rect 10599 11159 10625 11185
rect 10625 11159 10626 11185
rect 10598 11158 10626 11159
rect 10766 11158 10794 11186
rect 10486 11102 10514 11130
rect 9758 10934 9786 10962
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10486 10934 10514 10962
rect 10710 10934 10738 10962
rect 10374 10878 10402 10906
rect 9534 10038 9562 10066
rect 9590 10009 9618 10010
rect 9590 9983 9591 10009
rect 9591 9983 9617 10009
rect 9617 9983 9618 10009
rect 9590 9982 9618 9983
rect 9478 9870 9506 9898
rect 9422 9142 9450 9170
rect 9534 9030 9562 9058
rect 9366 8833 9394 8834
rect 9366 8807 9367 8833
rect 9367 8807 9393 8833
rect 9393 8807 9394 8833
rect 9366 8806 9394 8807
rect 9590 9310 9618 9338
rect 9310 8638 9338 8666
rect 9254 8441 9282 8442
rect 9254 8415 9255 8441
rect 9255 8415 9281 8441
rect 9281 8415 9282 8441
rect 9254 8414 9282 8415
rect 8862 7993 8890 7994
rect 8862 7967 8863 7993
rect 8863 7967 8889 7993
rect 8889 7967 8890 7993
rect 8862 7966 8890 7967
rect 8750 7574 8778 7602
rect 9646 8974 9674 9002
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9814 9673 9842 9674
rect 9814 9647 9815 9673
rect 9815 9647 9841 9673
rect 9841 9647 9842 9673
rect 9814 9646 9842 9647
rect 9870 10094 9898 10122
rect 10094 10094 10122 10122
rect 10150 9982 10178 10010
rect 10206 10094 10234 10122
rect 9926 9814 9954 9842
rect 10094 9758 10122 9786
rect 9926 9646 9954 9674
rect 10038 9702 10066 9730
rect 10430 10262 10458 10290
rect 10766 10094 10794 10122
rect 10934 11241 10962 11242
rect 10934 11215 10935 11241
rect 10935 11215 10961 11241
rect 10961 11215 10962 11241
rect 10934 11214 10962 11215
rect 11046 11214 11074 11242
rect 10038 9534 10066 9562
rect 10206 9561 10234 9562
rect 10206 9535 10207 9561
rect 10207 9535 10233 9561
rect 10233 9535 10234 9561
rect 10206 9534 10234 9535
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9758 9310 9786 9338
rect 9870 9225 9898 9226
rect 9870 9199 9871 9225
rect 9871 9199 9897 9225
rect 9897 9199 9898 9225
rect 9870 9198 9898 9199
rect 9702 8806 9730 8834
rect 10094 9225 10122 9226
rect 10094 9199 10095 9225
rect 10095 9199 10121 9225
rect 10121 9199 10122 9225
rect 10094 9198 10122 9199
rect 10878 9870 10906 9898
rect 10654 9142 10682 9170
rect 10374 9086 10402 9114
rect 10206 9030 10234 9058
rect 10150 8918 10178 8946
rect 10766 9030 10794 9058
rect 10766 8833 10794 8834
rect 10766 8807 10767 8833
rect 10767 8807 10793 8833
rect 10793 8807 10794 8833
rect 10766 8806 10794 8807
rect 11158 11550 11186 11578
rect 11158 10990 11186 11018
rect 11102 10934 11130 10962
rect 11662 12473 11690 12474
rect 11662 12447 11663 12473
rect 11663 12447 11689 12473
rect 11689 12447 11690 12473
rect 11662 12446 11690 12447
rect 11774 11633 11802 11634
rect 11774 11607 11775 11633
rect 11775 11607 11801 11633
rect 11801 11607 11802 11633
rect 11774 11606 11802 11607
rect 11942 13006 11970 13034
rect 13006 13873 13034 13874
rect 13006 13847 13007 13873
rect 13007 13847 13033 13873
rect 13033 13847 13034 13873
rect 13006 13846 13034 13847
rect 12726 13790 12754 13818
rect 12390 13537 12418 13538
rect 12390 13511 12391 13537
rect 12391 13511 12417 13537
rect 12417 13511 12418 13537
rect 12390 13510 12418 13511
rect 12334 13286 12362 13314
rect 14574 18745 14602 18746
rect 14574 18719 14575 18745
rect 14575 18719 14601 18745
rect 14601 18719 14602 18745
rect 14574 18718 14602 18719
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 13174 13510 13202 13538
rect 13118 13398 13146 13426
rect 12894 13286 12922 13314
rect 12614 13145 12642 13146
rect 12614 13119 12615 13145
rect 12615 13119 12641 13145
rect 12641 13119 12642 13145
rect 12614 13118 12642 13119
rect 12390 12697 12418 12698
rect 12390 12671 12391 12697
rect 12391 12671 12417 12697
rect 12417 12671 12418 12697
rect 12390 12670 12418 12671
rect 12950 13145 12978 13146
rect 12950 13119 12951 13145
rect 12951 13119 12977 13145
rect 12977 13119 12978 13145
rect 12950 13118 12978 13119
rect 12894 11942 12922 11970
rect 12166 11633 12194 11634
rect 12166 11607 12167 11633
rect 12167 11607 12193 11633
rect 12193 11607 12194 11633
rect 12166 11606 12194 11607
rect 12670 11830 12698 11858
rect 11382 11241 11410 11242
rect 11382 11215 11383 11241
rect 11383 11215 11409 11241
rect 11409 11215 11410 11241
rect 11382 11214 11410 11215
rect 11214 10822 11242 10850
rect 11326 10793 11354 10794
rect 11326 10767 11327 10793
rect 11327 10767 11353 10793
rect 11353 10767 11354 10793
rect 11326 10766 11354 10767
rect 11214 10009 11242 10010
rect 11214 9983 11215 10009
rect 11215 9983 11241 10009
rect 11241 9983 11242 10009
rect 11214 9982 11242 9983
rect 11662 11214 11690 11242
rect 11494 11129 11522 11130
rect 11494 11103 11495 11129
rect 11495 11103 11521 11129
rect 11521 11103 11522 11129
rect 11494 11102 11522 11103
rect 11774 10878 11802 10906
rect 11550 10822 11578 10850
rect 11774 10710 11802 10738
rect 11046 9534 11074 9562
rect 11046 9113 11074 9114
rect 11046 9087 11047 9113
rect 11047 9087 11073 9113
rect 11073 9087 11074 9113
rect 11046 9086 11074 9087
rect 10878 8918 10906 8946
rect 11158 9086 11186 9114
rect 11214 9030 11242 9058
rect 9926 8721 9954 8722
rect 9926 8695 9927 8721
rect 9927 8695 9953 8721
rect 9953 8695 9954 8721
rect 9926 8694 9954 8695
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 11270 8638 11298 8666
rect 11550 10598 11578 10626
rect 11886 10598 11914 10626
rect 11774 10318 11802 10346
rect 12166 11158 12194 11186
rect 12782 11718 12810 11746
rect 13286 13286 13314 13314
rect 13230 13257 13258 13258
rect 13230 13231 13231 13257
rect 13231 13231 13257 13257
rect 13257 13231 13258 13257
rect 13230 13230 13258 13231
rect 14014 13537 14042 13538
rect 14014 13511 14015 13537
rect 14015 13511 14041 13537
rect 14041 13511 14042 13537
rect 14014 13510 14042 13511
rect 13566 13286 13594 13314
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 14294 13510 14322 13538
rect 14910 13510 14938 13538
rect 14070 13230 14098 13258
rect 13398 13145 13426 13146
rect 13398 13119 13399 13145
rect 13399 13119 13425 13145
rect 13425 13119 13426 13145
rect 13398 13118 13426 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 13902 12278 13930 12306
rect 13790 11969 13818 11970
rect 13790 11943 13791 11969
rect 13791 11943 13817 11969
rect 13817 11943 13818 11969
rect 13790 11942 13818 11943
rect 14686 12305 14714 12306
rect 14686 12279 14687 12305
rect 14687 12279 14713 12305
rect 14713 12279 14714 12305
rect 14686 12278 14714 12279
rect 13174 11718 13202 11746
rect 13062 11606 13090 11634
rect 12166 11073 12194 11074
rect 12166 11047 12167 11073
rect 12167 11047 12193 11073
rect 12193 11047 12194 11073
rect 12166 11046 12194 11047
rect 11998 10990 12026 11018
rect 12054 10822 12082 10850
rect 12166 10318 12194 10346
rect 11774 9646 11802 9674
rect 11662 9422 11690 9450
rect 11382 9086 11410 9114
rect 11606 9142 11634 9170
rect 11830 9310 11858 9338
rect 11550 8974 11578 9002
rect 11718 9030 11746 9058
rect 11662 8833 11690 8834
rect 11662 8807 11663 8833
rect 11663 8807 11689 8833
rect 11689 8807 11690 8833
rect 11662 8806 11690 8807
rect 9254 7574 9282 7602
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10318 7574 10346 7602
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 8750 1806 8778 1834
rect 10486 7574 10514 7602
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10094 6817 10122 6818
rect 10094 6791 10095 6817
rect 10095 6791 10121 6817
rect 10121 6791 10122 6817
rect 10094 6790 10122 6791
rect 10710 6790 10738 6818
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9758 2030 9786 2058
rect 9310 1833 9338 1834
rect 9310 1807 9311 1833
rect 9311 1807 9337 1833
rect 9337 1807 9338 1833
rect 9310 1806 9338 1807
rect 10374 2057 10402 2058
rect 10374 2031 10375 2057
rect 10375 2031 10401 2057
rect 10401 2031 10402 2057
rect 10374 2030 10402 2031
rect 11606 8638 11634 8666
rect 12054 9646 12082 9674
rect 12110 9870 12138 9898
rect 12110 9534 12138 9562
rect 12222 10065 12250 10066
rect 12222 10039 12223 10065
rect 12223 10039 12249 10065
rect 12249 10039 12250 10065
rect 12222 10038 12250 10039
rect 12614 10793 12642 10794
rect 12614 10767 12615 10793
rect 12615 10767 12641 10793
rect 12641 10767 12642 10793
rect 12614 10766 12642 10767
rect 12670 10038 12698 10066
rect 12950 11185 12978 11186
rect 12950 11159 12951 11185
rect 12951 11159 12977 11185
rect 12977 11159 12978 11185
rect 12950 11158 12978 11159
rect 13062 11129 13090 11130
rect 13062 11103 13063 11129
rect 13063 11103 13089 11129
rect 13089 11103 13090 11129
rect 13062 11102 13090 11103
rect 12726 11046 12754 11074
rect 12334 9982 12362 10010
rect 12222 9617 12250 9618
rect 12222 9591 12223 9617
rect 12223 9591 12249 9617
rect 12249 9591 12250 9617
rect 12222 9590 12250 9591
rect 12502 9534 12530 9562
rect 12110 9169 12138 9170
rect 12110 9143 12111 9169
rect 12111 9143 12137 9169
rect 12137 9143 12138 9169
rect 12110 9142 12138 9143
rect 12054 9086 12082 9114
rect 11942 8974 11970 9002
rect 12166 8497 12194 8498
rect 12166 8471 12167 8497
rect 12167 8471 12193 8497
rect 12193 8471 12194 8497
rect 12166 8470 12194 8471
rect 11718 8385 11746 8386
rect 11718 8359 11719 8385
rect 11719 8359 11745 8385
rect 11745 8359 11746 8385
rect 11718 8358 11746 8359
rect 12278 9086 12306 9114
rect 12334 9030 12362 9058
rect 12838 10990 12866 11018
rect 12838 10150 12866 10178
rect 13454 11857 13482 11858
rect 13454 11831 13455 11857
rect 13455 11831 13481 11857
rect 13481 11831 13482 11857
rect 13454 11830 13482 11831
rect 14406 11689 14434 11690
rect 14406 11663 14407 11689
rect 14407 11663 14433 11689
rect 14433 11663 14434 11689
rect 14406 11662 14434 11663
rect 13734 11606 13762 11634
rect 13398 11241 13426 11242
rect 13398 11215 13399 11241
rect 13399 11215 13425 11241
rect 13425 11215 13426 11241
rect 13398 11214 13426 11215
rect 13342 10710 13370 10738
rect 13398 10345 13426 10346
rect 13398 10319 13399 10345
rect 13399 10319 13425 10345
rect 13425 10319 13426 10345
rect 13398 10318 13426 10319
rect 13622 10598 13650 10626
rect 13902 11550 13930 11578
rect 14182 11550 14210 11578
rect 14014 11129 14042 11130
rect 14014 11103 14015 11129
rect 14015 11103 14041 11129
rect 14041 11103 14042 11129
rect 14014 11102 14042 11103
rect 20006 12446 20034 12474
rect 18830 12278 18858 12306
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 14910 11662 14938 11690
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 13734 10374 13762 10402
rect 13790 10766 13818 10794
rect 13566 10345 13594 10346
rect 13566 10319 13567 10345
rect 13567 10319 13593 10345
rect 13593 10319 13594 10345
rect 13566 10318 13594 10319
rect 14294 10766 14322 10794
rect 13902 10598 13930 10626
rect 13846 10401 13874 10402
rect 13846 10375 13847 10401
rect 13847 10375 13873 10401
rect 13873 10375 13874 10401
rect 13846 10374 13874 10375
rect 13510 10289 13538 10290
rect 13510 10263 13511 10289
rect 13511 10263 13537 10289
rect 13537 10263 13538 10289
rect 13510 10262 13538 10263
rect 13286 10038 13314 10066
rect 13230 9617 13258 9618
rect 13230 9591 13231 9617
rect 13231 9591 13257 9617
rect 13257 9591 13258 9617
rect 13230 9590 13258 9591
rect 13342 9590 13370 9618
rect 12726 9422 12754 9450
rect 12614 9225 12642 9226
rect 12614 9199 12615 9225
rect 12615 9199 12641 9225
rect 12641 9199 12642 9225
rect 12614 9198 12642 9199
rect 12670 9113 12698 9114
rect 12670 9087 12671 9113
rect 12671 9087 12697 9113
rect 12697 9087 12698 9113
rect 12670 9086 12698 9087
rect 13342 9422 13370 9450
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 20006 10430 20034 10458
rect 13510 9617 13538 9618
rect 13510 9591 13511 9617
rect 13511 9591 13537 9617
rect 13537 9591 13538 9617
rect 13510 9590 13538 9591
rect 13118 9030 13146 9058
rect 13174 9142 13202 9170
rect 12614 8777 12642 8778
rect 12614 8751 12615 8777
rect 12615 8751 12641 8777
rect 12641 8751 12642 8777
rect 12614 8750 12642 8751
rect 12222 8134 12250 8162
rect 12558 8358 12586 8386
rect 12166 8049 12194 8050
rect 12166 8023 12167 8049
rect 12167 8023 12193 8049
rect 12193 8023 12194 8049
rect 12166 8022 12194 8023
rect 11662 7574 11690 7602
rect 11886 7601 11914 7602
rect 11886 7575 11887 7601
rect 11887 7575 11913 7601
rect 11913 7575 11914 7601
rect 11886 7574 11914 7575
rect 11494 7518 11522 7546
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 13398 9086 13426 9114
rect 13342 8862 13370 8890
rect 13230 8777 13258 8778
rect 13230 8751 13231 8777
rect 13231 8751 13257 8777
rect 13257 8751 13258 8777
rect 13230 8750 13258 8751
rect 12782 8441 12810 8442
rect 12782 8415 12783 8441
rect 12783 8415 12809 8441
rect 12809 8415 12810 8441
rect 12782 8414 12810 8415
rect 12782 8022 12810 8050
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14294 8889 14322 8890
rect 14294 8863 14295 8889
rect 14295 8863 14321 8889
rect 14321 8863 14322 8889
rect 14294 8862 14322 8863
rect 14294 8694 14322 8722
rect 13622 8470 13650 8498
rect 18830 8694 18858 8722
rect 14126 8414 14154 8442
rect 13958 8358 13986 8386
rect 13846 8161 13874 8162
rect 13846 8135 13847 8161
rect 13847 8135 13873 8161
rect 13873 8135 13874 8161
rect 13846 8134 13874 8135
rect 13622 8105 13650 8106
rect 13622 8079 13623 8105
rect 13623 8079 13649 8105
rect 13649 8079 13650 8105
rect 13622 8078 13650 8079
rect 13398 8022 13426 8050
rect 11494 6902 11522 6930
rect 11774 6929 11802 6930
rect 11774 6903 11775 6929
rect 11775 6903 11801 6929
rect 11801 6903 11802 6929
rect 11774 6902 11802 6903
rect 11382 6790 11410 6818
rect 13790 8049 13818 8050
rect 13790 8023 13791 8049
rect 13791 8023 13817 8049
rect 13817 8023 13818 8049
rect 13790 8022 13818 8023
rect 14238 8385 14266 8386
rect 14238 8359 14239 8385
rect 14239 8359 14265 8385
rect 14265 8359 14266 8385
rect 14238 8358 14266 8359
rect 20006 8750 20034 8778
rect 18886 8358 18914 8386
rect 20006 8414 20034 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 18830 8078 18858 8106
rect 20006 8105 20034 8106
rect 20006 8079 20007 8105
rect 20007 8079 20033 8105
rect 20033 8079 20034 8105
rect 20006 8078 20034 8079
rect 12222 7574 12250 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 11774 2590 11802 2618
rect 11438 1806 11466 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12390 2617 12418 2618
rect 12390 2591 12391 2617
rect 12391 2591 12417 2617
rect 12417 2591 12418 2617
rect 12390 2590 12418 2591
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 10761 19110 10766 19138
rect 10794 19110 11214 19138
rect 11242 19110 11247 19138
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 13449 19110 13454 19138
rect 13482 19110 14686 19138
rect 14714 19110 14719 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 12441 18718 12446 18746
rect 12474 18718 13118 18746
rect 13146 18718 13151 18746
rect 13785 18718 13790 18746
rect 13818 18718 14574 18746
rect 14602 18718 14607 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 0 18186 400 18200
rect 0 18158 854 18186
rect 882 18158 887 18186
rect 0 18144 400 18158
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 10817 14238 10822 14266
rect 10850 14238 12614 14266
rect 12642 14238 12782 14266
rect 12810 14238 12815 14266
rect 0 14154 400 14168
rect 0 14126 2086 14154
rect 2114 14126 2119 14154
rect 0 14112 400 14126
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2137 13902 2142 13930
rect 2170 13902 7630 13930
rect 7658 13902 7663 13930
rect 10649 13902 10654 13930
rect 10682 13902 11102 13930
rect 11130 13902 11135 13930
rect 11433 13902 11438 13930
rect 11466 13902 12166 13930
rect 12194 13902 12199 13930
rect 9361 13846 9366 13874
rect 9394 13846 10990 13874
rect 11018 13846 11023 13874
rect 12105 13846 12110 13874
rect 12138 13846 13006 13874
rect 13034 13846 13039 13874
rect 8913 13790 8918 13818
rect 8946 13790 11214 13818
rect 11242 13790 12054 13818
rect 12082 13790 12726 13818
rect 12754 13790 12759 13818
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 2137 13510 2142 13538
rect 2170 13510 7294 13538
rect 7322 13510 7327 13538
rect 12385 13510 12390 13538
rect 12418 13510 13174 13538
rect 13202 13510 14014 13538
rect 14042 13510 14294 13538
rect 14322 13510 14910 13538
rect 14938 13510 14943 13538
rect 0 13482 400 13496
rect 0 13454 966 13482
rect 994 13454 999 13482
rect 0 13440 400 13454
rect 11937 13398 11942 13426
rect 11970 13398 13118 13426
rect 13146 13398 13151 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 12329 13286 12334 13314
rect 12362 13286 12894 13314
rect 12922 13286 13286 13314
rect 13314 13286 13566 13314
rect 13594 13286 13599 13314
rect 10593 13230 10598 13258
rect 10626 13230 10878 13258
rect 10906 13230 10911 13258
rect 13225 13230 13230 13258
rect 13258 13230 14070 13258
rect 14098 13230 14103 13258
rect 0 13146 400 13160
rect 0 13118 1022 13146
rect 1050 13118 1055 13146
rect 2137 13118 2142 13146
rect 2170 13118 5950 13146
rect 5978 13118 7462 13146
rect 7490 13118 7742 13146
rect 7770 13118 7775 13146
rect 8689 13118 8694 13146
rect 8722 13118 9142 13146
rect 9170 13118 10598 13146
rect 10626 13118 10631 13146
rect 11881 13118 11886 13146
rect 11914 13118 12614 13146
rect 12642 13118 12647 13146
rect 12945 13118 12950 13146
rect 12978 13118 13398 13146
rect 13426 13118 13431 13146
rect 0 13104 400 13118
rect 7401 13062 7406 13090
rect 7434 13062 7630 13090
rect 7658 13062 8022 13090
rect 8050 13062 9366 13090
rect 9394 13062 9399 13090
rect 9025 13006 9030 13034
rect 9058 13006 9198 13034
rect 9226 13006 9231 13034
rect 9305 13006 9310 13034
rect 9338 13006 9534 13034
rect 9562 13006 11942 13034
rect 11970 13006 11975 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 0 12810 400 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 7961 12782 7966 12810
rect 7994 12782 8750 12810
rect 8778 12782 8783 12810
rect 10593 12782 10598 12810
rect 10626 12782 11830 12810
rect 11858 12782 11863 12810
rect 0 12768 400 12782
rect 10369 12726 10374 12754
rect 10402 12726 11158 12754
rect 11186 12726 11662 12754
rect 11690 12726 11695 12754
rect 10201 12670 10206 12698
rect 10234 12670 11270 12698
rect 11298 12670 12390 12698
rect 12418 12670 12423 12698
rect 10145 12614 10150 12642
rect 10178 12614 10710 12642
rect 10738 12614 10743 12642
rect 10201 12558 10206 12586
rect 10234 12558 10239 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 7793 12502 7798 12530
rect 7826 12502 8806 12530
rect 8834 12502 9646 12530
rect 9674 12502 9679 12530
rect 10206 12474 10234 12558
rect 20600 12474 21000 12488
rect 6953 12446 6958 12474
rect 6986 12446 7742 12474
rect 7770 12446 7775 12474
rect 7905 12446 7910 12474
rect 7938 12446 9086 12474
rect 9114 12446 9119 12474
rect 9865 12446 9870 12474
rect 9898 12446 10234 12474
rect 10985 12446 10990 12474
rect 11018 12446 11662 12474
rect 11690 12446 11695 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 20600 12432 21000 12446
rect 13897 12278 13902 12306
rect 13930 12278 14686 12306
rect 14714 12278 18830 12306
rect 18858 12278 18863 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 2137 11942 2142 11970
rect 2170 11942 5558 11970
rect 5586 11942 6846 11970
rect 6874 11942 6879 11970
rect 12889 11942 12894 11970
rect 12922 11942 13790 11970
rect 13818 11942 13823 11970
rect 6897 11886 6902 11914
rect 6930 11886 7742 11914
rect 7770 11886 7775 11914
rect 7233 11830 7238 11858
rect 7266 11830 8022 11858
rect 8050 11830 8055 11858
rect 12665 11830 12670 11858
rect 12698 11830 13454 11858
rect 13482 11830 13487 11858
rect 0 11802 400 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 12777 11718 12782 11746
rect 12810 11718 13174 11746
rect 13202 11718 13207 11746
rect 6617 11662 6622 11690
rect 6650 11662 8078 11690
rect 8106 11662 8111 11690
rect 8185 11662 8190 11690
rect 8218 11662 8638 11690
rect 8666 11662 8671 11690
rect 8745 11662 8750 11690
rect 8778 11662 9310 11690
rect 9338 11662 9343 11690
rect 10425 11662 10430 11690
rect 10458 11662 10710 11690
rect 10738 11662 10743 11690
rect 14401 11662 14406 11690
rect 14434 11662 14910 11690
rect 14938 11662 14943 11690
rect 8078 11634 8106 11662
rect 8078 11606 9870 11634
rect 9898 11606 9903 11634
rect 11769 11606 11774 11634
rect 11802 11606 12166 11634
rect 12194 11606 12199 11634
rect 13057 11606 13062 11634
rect 13090 11606 13734 11634
rect 13762 11606 13767 11634
rect 10705 11550 10710 11578
rect 10738 11550 11158 11578
rect 11186 11550 11191 11578
rect 13897 11550 13902 11578
rect 13930 11550 14182 11578
rect 14210 11550 18830 11578
rect 18858 11550 18863 11578
rect 20600 11466 21000 11480
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9753 11214 9758 11242
rect 9786 11214 10934 11242
rect 10962 11214 10967 11242
rect 11041 11214 11046 11242
rect 11074 11214 11382 11242
rect 11410 11214 11662 11242
rect 11690 11214 13398 11242
rect 13426 11214 13431 11242
rect 8297 11158 8302 11186
rect 8330 11158 9086 11186
rect 9114 11158 9119 11186
rect 9305 11158 9310 11186
rect 9338 11158 9814 11186
rect 9842 11158 9847 11186
rect 10066 11158 10598 11186
rect 10626 11158 10631 11186
rect 10761 11158 10766 11186
rect 10794 11158 10799 11186
rect 12161 11158 12166 11186
rect 12194 11158 12950 11186
rect 12978 11158 12983 11186
rect 10066 11130 10094 11158
rect 10766 11130 10794 11158
rect 9865 11102 9870 11130
rect 9898 11102 10094 11130
rect 10481 11102 10486 11130
rect 10514 11102 11494 11130
rect 11522 11102 11527 11130
rect 13057 11102 13062 11130
rect 13090 11102 14014 11130
rect 14042 11102 14047 11130
rect 10033 11046 10038 11074
rect 10066 11046 10402 11074
rect 12161 11046 12166 11074
rect 12194 11046 12726 11074
rect 12754 11046 12759 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 9417 10934 9422 10962
rect 9450 10934 9758 10962
rect 9786 10934 9791 10962
rect 10374 10906 10402 11046
rect 11153 10990 11158 11018
rect 11186 10990 11998 11018
rect 12026 10990 12838 11018
rect 12866 10990 12871 11018
rect 10481 10934 10486 10962
rect 10514 10934 10710 10962
rect 10738 10934 11102 10962
rect 11130 10934 13566 10962
rect 13594 10934 13599 10962
rect 6561 10878 6566 10906
rect 6594 10878 6902 10906
rect 6930 10878 6935 10906
rect 8409 10878 8414 10906
rect 8442 10878 9590 10906
rect 9618 10878 9623 10906
rect 10369 10878 10374 10906
rect 10402 10878 11774 10906
rect 11802 10878 11807 10906
rect 8465 10822 8470 10850
rect 8498 10822 8806 10850
rect 8834 10822 9142 10850
rect 9170 10822 9175 10850
rect 11209 10822 11214 10850
rect 11242 10822 11550 10850
rect 11578 10822 12054 10850
rect 12082 10822 12087 10850
rect 2137 10766 2142 10794
rect 2170 10766 4998 10794
rect 5026 10766 5031 10794
rect 8297 10766 8302 10794
rect 8330 10766 8750 10794
rect 8778 10766 8783 10794
rect 11321 10766 11326 10794
rect 11354 10766 12614 10794
rect 12642 10766 12647 10794
rect 13785 10766 13790 10794
rect 13818 10766 14294 10794
rect 14322 10766 18830 10794
rect 18858 10766 18863 10794
rect 11769 10710 11774 10738
rect 11802 10710 13342 10738
rect 13370 10710 13375 10738
rect 11545 10598 11550 10626
rect 11578 10598 11886 10626
rect 11914 10598 13622 10626
rect 13650 10598 13902 10626
rect 13930 10598 13935 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7905 10486 7910 10514
rect 7938 10486 8582 10514
rect 8610 10486 10094 10514
rect 0 10458 400 10472
rect 0 10430 966 10458
rect 994 10430 999 10458
rect 4993 10430 4998 10458
rect 5026 10430 6678 10458
rect 6706 10430 6711 10458
rect 0 10416 400 10430
rect 10066 10402 10094 10486
rect 20600 10458 21000 10472
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 20600 10416 21000 10430
rect 7961 10374 7966 10402
rect 7994 10374 8582 10402
rect 8610 10374 9086 10402
rect 9114 10374 9119 10402
rect 10066 10374 13734 10402
rect 13762 10374 13846 10402
rect 13874 10374 13879 10402
rect 9305 10318 9310 10346
rect 9338 10318 11774 10346
rect 11802 10318 11807 10346
rect 12161 10318 12166 10346
rect 12194 10318 13398 10346
rect 13426 10318 13431 10346
rect 13547 10318 13566 10346
rect 13594 10318 13599 10346
rect 2081 10262 2086 10290
rect 2114 10262 10430 10290
rect 10458 10262 10463 10290
rect 13426 10262 13510 10290
rect 13538 10262 13543 10290
rect 7793 10206 7798 10234
rect 7826 10206 8694 10234
rect 8722 10206 9310 10234
rect 9338 10206 9343 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 13426 10178 13454 10262
rect 12833 10150 12838 10178
rect 12866 10150 13454 10178
rect 7737 10094 7742 10122
rect 7770 10094 8246 10122
rect 8274 10094 8279 10122
rect 8745 10094 8750 10122
rect 8778 10094 9254 10122
rect 9282 10094 9870 10122
rect 9898 10094 9903 10122
rect 10089 10094 10094 10122
rect 10122 10094 10206 10122
rect 10234 10094 10766 10122
rect 10794 10094 10799 10122
rect 6393 10038 6398 10066
rect 6426 10038 7182 10066
rect 7210 10038 7215 10066
rect 8073 10038 8078 10066
rect 8106 10038 8862 10066
rect 8890 10038 9142 10066
rect 9170 10038 9175 10066
rect 9529 10038 9534 10066
rect 9562 10038 9730 10066
rect 12217 10038 12222 10066
rect 12250 10038 12670 10066
rect 12698 10038 13286 10066
rect 13314 10038 13319 10066
rect 7233 9982 7238 10010
rect 7266 9982 7574 10010
rect 7602 9982 7607 10010
rect 7905 9982 7910 10010
rect 7938 9982 8190 10010
rect 8218 9982 8806 10010
rect 8834 9982 8839 10010
rect 8969 9982 8974 10010
rect 9002 9982 9590 10010
rect 9618 9982 9623 10010
rect 8974 9954 9002 9982
rect 8241 9926 8246 9954
rect 8274 9926 9002 9954
rect 9137 9870 9142 9898
rect 9170 9870 9478 9898
rect 9506 9870 9511 9898
rect 9702 9842 9730 10038
rect 10145 9982 10150 10010
rect 10178 9982 11214 10010
rect 11242 9982 12334 10010
rect 12362 9982 12367 10010
rect 10873 9870 10878 9898
rect 10906 9870 12110 9898
rect 12138 9870 12143 9898
rect 9361 9814 9366 9842
rect 9394 9814 9926 9842
rect 9954 9814 9959 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 7177 9758 7182 9786
rect 7210 9758 10094 9786
rect 10122 9758 10127 9786
rect 10878 9730 10906 9870
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 10033 9702 10038 9730
rect 10066 9702 10906 9730
rect 9809 9646 9814 9674
rect 9842 9646 9847 9674
rect 9921 9646 9926 9674
rect 9954 9646 11774 9674
rect 11802 9646 12054 9674
rect 12082 9646 12087 9674
rect 9814 9618 9842 9646
rect 9814 9590 12222 9618
rect 12250 9590 13230 9618
rect 13258 9590 13263 9618
rect 13337 9590 13342 9618
rect 13370 9590 13510 9618
rect 13538 9590 13543 9618
rect 9193 9534 9198 9562
rect 9226 9534 10038 9562
rect 10066 9534 10071 9562
rect 10201 9534 10206 9562
rect 10234 9534 11046 9562
rect 11074 9534 11079 9562
rect 12105 9534 12110 9562
rect 12138 9534 12502 9562
rect 12530 9534 12535 9562
rect 11657 9422 11662 9450
rect 11690 9422 12726 9450
rect 12754 9422 13342 9450
rect 13370 9422 13375 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 8409 9310 8414 9338
rect 8442 9310 8918 9338
rect 8946 9310 9590 9338
rect 9618 9310 9758 9338
rect 9786 9310 11830 9338
rect 11858 9310 11863 9338
rect 6729 9254 6734 9282
rect 6762 9254 7182 9282
rect 7210 9254 7215 9282
rect 2137 9198 2142 9226
rect 2170 9198 5446 9226
rect 5474 9198 7126 9226
rect 7154 9198 7159 9226
rect 8409 9198 8414 9226
rect 8442 9198 8750 9226
rect 8778 9198 8974 9226
rect 9002 9198 9870 9226
rect 9898 9198 9903 9226
rect 10089 9198 10094 9226
rect 10122 9198 12614 9226
rect 12642 9198 12647 9226
rect 6897 9142 6902 9170
rect 6930 9142 7406 9170
rect 7434 9142 7439 9170
rect 9417 9142 9422 9170
rect 9450 9142 10570 9170
rect 10649 9142 10654 9170
rect 10682 9142 11606 9170
rect 11634 9142 11639 9170
rect 12105 9142 12110 9170
rect 12138 9142 13174 9170
rect 13202 9142 13207 9170
rect 0 9114 400 9128
rect 10542 9114 10570 9142
rect 0 9086 966 9114
rect 994 9086 999 9114
rect 9137 9086 9142 9114
rect 9170 9086 10374 9114
rect 10402 9086 10514 9114
rect 10542 9086 11046 9114
rect 11074 9086 11158 9114
rect 11186 9086 11382 9114
rect 11410 9086 11415 9114
rect 11494 9086 12054 9114
rect 12082 9086 12087 9114
rect 12273 9086 12278 9114
rect 12306 9086 12670 9114
rect 12698 9086 13398 9114
rect 13426 9086 13431 9114
rect 0 9072 400 9086
rect 10486 9058 10514 9086
rect 11494 9058 11522 9086
rect 9529 9030 9534 9058
rect 9562 9030 10206 9058
rect 10234 9030 10239 9058
rect 10486 9030 10766 9058
rect 10794 9030 10799 9058
rect 11209 9030 11214 9058
rect 11242 9030 11522 9058
rect 11713 9030 11718 9058
rect 11746 9030 12334 9058
rect 12362 9030 13118 9058
rect 13146 9030 13151 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9641 8974 9646 9002
rect 9674 8974 11550 9002
rect 11578 8974 11942 9002
rect 11970 8974 11975 9002
rect 10145 8918 10150 8946
rect 10178 8918 10878 8946
rect 10906 8918 10911 8946
rect 13337 8862 13342 8890
rect 13370 8862 14294 8890
rect 14322 8862 14327 8890
rect 2137 8806 2142 8834
rect 2170 8806 6342 8834
rect 6370 8806 8134 8834
rect 8162 8806 8167 8834
rect 8241 8806 8246 8834
rect 8274 8806 9198 8834
rect 9226 8806 9231 8834
rect 9361 8806 9366 8834
rect 9394 8806 9702 8834
rect 9730 8806 9735 8834
rect 10761 8806 10766 8834
rect 10794 8806 11662 8834
rect 11690 8806 11695 8834
rect 9366 8778 9394 8806
rect 20600 8778 21000 8792
rect 7233 8750 7238 8778
rect 7266 8750 8078 8778
rect 8106 8750 8111 8778
rect 8297 8750 8302 8778
rect 8330 8750 8694 8778
rect 8722 8750 8727 8778
rect 9137 8750 9142 8778
rect 9170 8750 9394 8778
rect 12609 8750 12614 8778
rect 12642 8750 13230 8778
rect 13258 8750 13263 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 6841 8694 6846 8722
rect 6874 8694 8918 8722
rect 8946 8694 8951 8722
rect 9193 8694 9198 8722
rect 9226 8694 9926 8722
rect 9954 8694 9959 8722
rect 14289 8694 14294 8722
rect 14322 8694 18830 8722
rect 18858 8694 18863 8722
rect 9198 8638 9310 8666
rect 9338 8638 9343 8666
rect 11265 8638 11270 8666
rect 11298 8638 11606 8666
rect 11634 8638 11639 8666
rect 9198 8610 9226 8638
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 9193 8582 9198 8610
rect 9226 8582 9231 8610
rect 12161 8470 12166 8498
rect 12194 8470 13622 8498
rect 13650 8470 13655 8498
rect 0 8442 400 8456
rect 20600 8442 21000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 7233 8414 7238 8442
rect 7266 8414 7462 8442
rect 7490 8414 7798 8442
rect 7826 8414 8022 8442
rect 8050 8414 9254 8442
rect 9282 8414 9287 8442
rect 12777 8414 12782 8442
rect 12810 8414 14126 8442
rect 14154 8414 14159 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 0 8400 400 8414
rect 20600 8400 21000 8414
rect 11713 8358 11718 8386
rect 11746 8358 12558 8386
rect 12586 8358 12591 8386
rect 13953 8358 13958 8386
rect 13986 8358 14238 8386
rect 14266 8358 18886 8386
rect 18914 8358 18919 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 12217 8134 12222 8162
rect 12250 8134 13846 8162
rect 13874 8134 13879 8162
rect 20600 8106 21000 8120
rect 13617 8078 13622 8106
rect 13650 8078 18830 8106
rect 18858 8078 18863 8106
rect 20001 8078 20006 8106
rect 20034 8078 21000 8106
rect 20600 8064 21000 8078
rect 12161 8022 12166 8050
rect 12194 8022 12782 8050
rect 12810 8022 12815 8050
rect 13393 8022 13398 8050
rect 13426 8022 13790 8050
rect 13818 8022 13823 8050
rect 7569 7966 7574 7994
rect 7602 7966 8862 7994
rect 8890 7966 8895 7994
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 8745 7574 8750 7602
rect 8778 7574 9254 7602
rect 9282 7574 10318 7602
rect 10346 7574 10351 7602
rect 10481 7574 10486 7602
rect 10514 7574 11522 7602
rect 11657 7574 11662 7602
rect 11690 7574 11886 7602
rect 11914 7574 12222 7602
rect 12250 7574 12255 7602
rect 11494 7546 11522 7574
rect 11489 7518 11494 7546
rect 11522 7518 11527 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 11489 6902 11494 6930
rect 11522 6902 11774 6930
rect 11802 6902 11807 6930
rect 10089 6790 10094 6818
rect 10122 6790 10710 6818
rect 10738 6790 11382 6818
rect 11410 6790 11415 6818
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 11769 2590 11774 2618
rect 11802 2590 12390 2618
rect 12418 2590 12423 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 9753 2030 9758 2058
rect 9786 2030 10374 2058
rect 10402 2030 10407 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 8745 1806 8750 1834
rect 8778 1806 9310 1834
rect 9338 1806 9343 1834
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 13566 10934 13594 10962
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 13566 10318 13594 10346
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 9904 10206 10064 10962
rect 13566 10962 13594 10967
rect 13566 10346 13594 10934
rect 13566 10313 13594 10318
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8176 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9184 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10024 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform -1 0 11312 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13664 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_
timestamp 1698175906
transform -1 0 12152 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _105_
timestamp 1698175906
transform -1 0 8176 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _106_
timestamp 1698175906
transform 1 0 9016 0 1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform -1 0 9016 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform -1 0 8512 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8680 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _111_
timestamp 1698175906
transform -1 0 10808 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11984 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _113_
timestamp 1698175906
transform -1 0 10248 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9128 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _116_
timestamp 1698175906
transform -1 0 12096 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9520 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13160 0 1 9408
box -43 -43 1891 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 12432 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _121_
timestamp 1698175906
transform 1 0 11312 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _122_
timestamp 1698175906
transform -1 0 11536 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10920 0 1 11760
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11536 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _126_
timestamp 1698175906
transform 1 0 9184 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _128_
timestamp 1698175906
transform 1 0 8176 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform -1 0 9576 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform -1 0 8904 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_
timestamp 1698175906
transform -1 0 8288 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 11424 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10416 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform -1 0 7840 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform -1 0 7336 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform -1 0 9408 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _137_
timestamp 1698175906
transform -1 0 9016 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform -1 0 8008 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _139_
timestamp 1698175906
transform 1 0 7504 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _140_
timestamp 1698175906
transform -1 0 7056 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform -1 0 6832 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform -1 0 6552 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10248 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _144_
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 13720 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform 1 0 11536 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _147_
timestamp 1698175906
transform 1 0 11872 0 -1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform 1 0 11984 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _149_
timestamp 1698175906
transform 1 0 13160 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _150_
timestamp 1698175906
transform 1 0 11984 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10024 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _153_
timestamp 1698175906
transform 1 0 10360 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 1107 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 1051 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _156_
timestamp 1698175906
transform -1 0 10248 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _157_
timestamp 1698175906
transform 1 0 11312 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _159_
timestamp 1698175906
transform 1 0 9520 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9520 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _161_
timestamp 1698175906
transform 1 0 11872 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform -1 0 11872 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _163_
timestamp 1698175906
transform 1 0 10976 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10696 0 1 8624
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1698175906
transform -1 0 11200 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 7000 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 6776 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform 1 0 13776 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13160 0 1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1698175906
transform -1 0 13160 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform 1 0 13720 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _172_
timestamp 1698175906
transform 1 0 13272 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _173_
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _174_
timestamp 1698175906
transform 1 0 12040 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698175906
transform -1 0 13384 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _176_
timestamp 1698175906
transform -1 0 12264 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 7280 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _178_
timestamp 1698175906
transform -1 0 10304 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _179_
timestamp 1698175906
transform -1 0 9296 0 1 8624
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform -1 0 6944 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform -1 0 12432 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _182_
timestamp 1698175906
transform 1 0 11032 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _183_
timestamp 1698175906
transform -1 0 12040 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform -1 0 13664 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _185_
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 9408 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _187_
timestamp 1698175906
transform -1 0 9128 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform -1 0 13496 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _189_
timestamp 1698175906
transform -1 0 12768 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7952 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_
timestamp 1698175906
transform 1 0 7168 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 13944 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _193_
timestamp 1698175906
transform -1 0 13776 0 1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform -1 0 11648 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform -1 0 14392 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 6776 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _200_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7560 0 -1 13328
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform 1 0 12712 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 12096 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 10360 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform -1 0 7112 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 13160 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform -1 0 7000 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 10696 0 1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 12264 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 7504 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 12768 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform -1 0 7896 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _220_
timestamp 1698175906
transform -1 0 12320 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _221_
timestamp 1698175906
transform -1 0 7896 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _222_
timestamp 1698175906
transform 1 0 12320 0 1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _223_
timestamp 1698175906
transform -1 0 7560 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 11760 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 14504 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 11648 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 8400 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 9128 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 8008 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 6552 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform -1 0 11032 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform -1 0 10360 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 14112 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 11984 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 7224 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 14392 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 14896 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 7392 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 12768 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 9240 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 14616 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 8008 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 14504 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 11424 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_158
timestamp 1698175906
transform 1 0 9520 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_162
timestamp 1698175906
transform 1 0 9744 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_189
timestamp 1698175906
transform 1 0 11256 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_205
timestamp 1698175906
transform 1 0 12152 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698175906
transform 1 0 11480 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_197
timestamp 1698175906
transform 1 0 11704 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_225
timestamp 1698175906
transform 1 0 13272 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_158 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_166
timestamp 1698175906
transform 1 0 9968 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_196
timestamp 1698175906
transform 1 0 11648 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_200
timestamp 1698175906
transform 1 0 11872 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 10360 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_193
timestamp 1698175906
transform 1 0 11480 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_201
timestamp 1698175906
transform 1 0 11928 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_204
timestamp 1698175906
transform 1 0 12096 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_236
timestamp 1698175906
transform 1 0 13888 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_171
timestamp 1698175906
transform 1 0 10248 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 12320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_220
timestamp 1698175906
transform 1 0 12992 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_229
timestamp 1698175906
transform 1 0 13496 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_261
timestamp 1698175906
transform 1 0 15288 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_164
timestamp 1698175906
transform 1 0 9856 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_193
timestamp 1698175906
transform 1 0 11480 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_201
timestamp 1698175906
transform 1 0 11928 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_203
timestamp 1698175906
transform 1 0 12040 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_238
timestamp 1698175906
transform 1 0 14000 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_96
timestamp 1698175906
transform 1 0 6048 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_129
timestamp 1698175906
transform 1 0 7896 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698175906
transform 1 0 8120 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 8344 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_151
timestamp 1698175906
transform 1 0 9128 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_155
timestamp 1698175906
transform 1 0 9352 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_171
timestamp 1698175906
transform 1 0 10248 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_179
timestamp 1698175906
transform 1 0 10696 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_181
timestamp 1698175906
transform 1 0 10808 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_214
timestamp 1698175906
transform 1 0 12656 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_244
timestamp 1698175906
transform 1 0 14336 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_248
timestamp 1698175906
transform 1 0 14560 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_112
timestamp 1698175906
transform 1 0 6944 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_120
timestamp 1698175906
transform 1 0 7392 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_128
timestamp 1698175906
transform 1 0 7840 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_140
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_144
timestamp 1698175906
transform 1 0 8736 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_146
timestamp 1698175906
transform 1 0 8848 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 10304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_205
timestamp 1698175906
transform 1 0 12152 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_207
timestamp 1698175906
transform 1 0 12264 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 14728 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 2240 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 4032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 4480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_118
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_122
timestamp 1698175906
transform 1 0 7504 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_130
timestamp 1698175906
transform 1 0 7952 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_153
timestamp 1698175906
transform 1 0 9240 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_161
timestamp 1698175906
transform 1 0 9688 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_171
timestamp 1698175906
transform 1 0 10248 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_179
timestamp 1698175906
transform 1 0 10696 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_183
timestamp 1698175906
transform 1 0 10920 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_198
timestamp 1698175906
transform 1 0 11760 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_245
timestamp 1698175906
transform 1 0 14392 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_249
timestamp 1698175906
transform 1 0 14616 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_265
timestamp 1698175906
transform 1 0 15512 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698175906
transform 1 0 15960 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 16184 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_139
timestamp 1698175906
transform 1 0 8456 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_183
timestamp 1698175906
transform 1 0 10920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_187
timestamp 1698175906
transform 1 0 11144 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_189
timestamp 1698175906
transform 1 0 11256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_231
timestamp 1698175906
transform 1 0 13608 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_239
timestamp 1698175906
transform 1 0 14056 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 14280 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_96
timestamp 1698175906
transform 1 0 6048 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_110
timestamp 1698175906
transform 1 0 6832 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_119
timestamp 1698175906
transform 1 0 7336 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_190
timestamp 1698175906
transform 1 0 11312 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_198
timestamp 1698175906
transform 1 0 11760 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 12320 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_245
timestamp 1698175906
transform 1 0 14392 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_249
timestamp 1698175906
transform 1 0 14616 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_265
timestamp 1698175906
transform 1 0 15512 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698175906
transform 1 0 15960 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 16184 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 16296 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_136
timestamp 1698175906
transform 1 0 8288 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_138
timestamp 1698175906
transform 1 0 8400 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_149
timestamp 1698175906
transform 1 0 9016 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_171
timestamp 1698175906
transform 1 0 10248 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_237
timestamp 1698175906
transform 1 0 13944 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 2240 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 4032 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 4480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698175906
transform 1 0 6496 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_107
timestamp 1698175906
transform 1 0 6664 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_123
timestamp 1698175906
transform 1 0 7560 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_127
timestamp 1698175906
transform 1 0 7784 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_262
timestamp 1698175906
transform 1 0 15344 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_123
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_131
timestamp 1698175906
transform 1 0 8008 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_135
timestamp 1698175906
transform 1 0 8232 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_137
timestamp 1698175906
transform 1 0 8344 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_140
timestamp 1698175906
transform 1 0 8512 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_210
timestamp 1698175906
transform 1 0 12432 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_239
timestamp 1698175906
transform 1 0 14056 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 8400 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_147
timestamp 1698175906
transform 1 0 8904 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_151
timestamp 1698175906
transform 1 0 9128 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_159
timestamp 1698175906
transform 1 0 9576 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_167
timestamp 1698175906
transform 1 0 10024 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_171
timestamp 1698175906
transform 1 0 10248 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_181
timestamp 1698175906
transform 1 0 10808 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_183
timestamp 1698175906
transform 1 0 10920 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_190
timestamp 1698175906
transform 1 0 11312 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_243
timestamp 1698175906
transform 1 0 14280 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_247
timestamp 1698175906
transform 1 0 14504 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_113
timestamp 1698175906
transform 1 0 7000 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_121
timestamp 1698175906
transform 1 0 7448 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_136
timestamp 1698175906
transform 1 0 8288 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698175906
transform 1 0 10080 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 10304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698175906
transform 1 0 10808 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_195
timestamp 1698175906
transform 1 0 11592 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_211
timestamp 1698175906
transform 1 0 12488 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_219
timestamp 1698175906
transform 1 0 12936 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_223
timestamp 1698175906
transform 1 0 13160 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698175906
transform 1 0 14000 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 14224 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 5152 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 5376 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_115
timestamp 1698175906
transform 1 0 7112 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_119
timestamp 1698175906
transform 1 0 7336 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_121
timestamp 1698175906
transform 1 0 7448 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_131
timestamp 1698175906
transform 1 0 8008 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_148
timestamp 1698175906
transform 1 0 8960 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_185
timestamp 1698175906
transform 1 0 11032 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_187
timestamp 1698175906
transform 1 0 11144 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_194
timestamp 1698175906
transform 1 0 11536 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_198
timestamp 1698175906
transform 1 0 11760 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 12208 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698175906
transform 1 0 12768 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_252
timestamp 1698175906
transform 1 0 14784 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_256
timestamp 1698175906
transform 1 0 15008 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_272
timestamp 1698175906
transform 1 0 15904 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698175906
transform 1 0 6776 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_114
timestamp 1698175906
transform 1 0 7056 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_151
timestamp 1698175906
transform 1 0 9128 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_155
timestamp 1698175906
transform 1 0 9352 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_163
timestamp 1698175906
transform 1 0 9800 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_211
timestamp 1698175906
transform 1 0 12488 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 14280 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_129
timestamp 1698175906
transform 1 0 7896 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698175906
transform 1 0 8120 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698175906
transform 1 0 8344 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_156
timestamp 1698175906
transform 1 0 9408 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_172
timestamp 1698175906
transform 1 0 10304 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_181
timestamp 1698175906
transform 1 0 10808 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_197
timestamp 1698175906
transform 1 0 11704 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698175906
transform 1 0 12152 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698175906
transform 1 0 12992 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_232
timestamp 1698175906
transform 1 0 13664 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_264
timestamp 1698175906
transform 1 0 15456 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 2240 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 2464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_115
timestamp 1698175906
transform 1 0 7112 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_155
timestamp 1698175906
transform 1 0 9352 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_163
timestamp 1698175906
transform 1 0 9800 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_193
timestamp 1698175906
transform 1 0 11480 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_197
timestamp 1698175906
transform 1 0 11704 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_236
timestamp 1698175906
transform 1 0 13888 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_240
timestamp 1698175906
transform 1 0 14112 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_28
timestamp 1698175906
transform 1 0 2240 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_60
timestamp 1698175906
transform 1 0 4032 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698175906
transform 1 0 4480 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_150
timestamp 1698175906
transform 1 0 9072 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_181
timestamp 1698175906
transform 1 0 10808 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_193
timestamp 1698175906
transform 1 0 11480 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_201
timestamp 1698175906
transform 1 0 11928 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_241
timestamp 1698175906
transform 1 0 14168 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_245
timestamp 1698175906
transform 1 0 14392 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_277
timestamp 1698175906
transform 1 0 16184 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 16296 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_214
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_218
timestamp 1698175906
transform 1 0 12880 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_234
timestamp 1698175906
transform 1 0 13776 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 14336 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 1008 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 1904 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 2352 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698175906
transform 1 0 12208 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_264
timestamp 1698175906
transform 1 0 15456 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_266
timestamp 1698175906
transform 1 0 15568 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698175906
transform 1 0 15792 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita47_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8512 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita47_26
timestamp 1698175906
transform -1 0 1008 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2240 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 14000 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 11816 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 -1 14112
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 9800 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 2240 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 2240 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 14112 400 14168 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 9072 400 9128 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 13776 20600 13832 21000 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 0 18144 400 18200 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 13440 20600 13496 21000 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 10416 400 10472 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 11172 14140 11172 14140 0 _000_
rlabel metal2 12684 13356 12684 13356 0 _001_
rlabel metal3 8372 12796 8372 12796 0 _002_
rlabel metal3 12936 8764 12936 8764 0 _003_
rlabel metal2 7420 8596 7420 8596 0 _004_
rlabel metal2 13328 9212 13328 9212 0 _005_
rlabel metal3 8232 7980 8232 7980 0 _006_
rlabel metal2 11172 7616 11172 7616 0 _007_
rlabel metal2 11900 10640 11900 10640 0 _008_
rlabel metal2 11284 12572 11284 12572 0 _009_
rlabel metal2 7252 11732 7252 11732 0 _010_
rlabel metal2 7084 10220 7084 10220 0 _011_
rlabel metal2 6916 12964 6916 12964 0 _012_
rlabel metal2 6300 10220 6300 10220 0 _013_
rlabel metal2 13188 8820 13188 8820 0 _014_
rlabel metal2 9996 13664 9996 13664 0 _015_
rlabel metal2 9100 7840 9100 7840 0 _016_
rlabel metal2 12572 8232 12572 8232 0 _017_
rlabel metal2 10836 8008 10836 8008 0 _018_
rlabel metal2 6524 11984 6524 11984 0 _019_
rlabel metal2 13020 11396 13020 11396 0 _020_
rlabel metal2 13636 12152 13636 12152 0 _021_
rlabel metal2 12124 13720 12124 13720 0 _022_
rlabel metal2 6692 8988 6692 8988 0 _023_
rlabel metal2 12684 11564 12684 11564 0 _024_
rlabel metal2 12348 9128 12348 9128 0 _025_
rlabel metal3 10780 12740 10780 12740 0 _026_
rlabel metal2 10808 11676 10808 11676 0 _027_
rlabel metal2 10556 13244 10556 13244 0 _028_
rlabel metal2 10668 13300 10668 13300 0 _029_
rlabel metal2 10164 13048 10164 13048 0 _030_
rlabel metal2 11452 9100 11452 9100 0 _031_
rlabel metal2 9380 8148 9380 8148 0 _032_
rlabel metal2 9436 8064 9436 8064 0 _033_
rlabel metal2 11956 8316 11956 8316 0 _034_
rlabel metal2 11004 8960 11004 8960 0 _035_
rlabel metal2 11032 8428 11032 8428 0 _036_
rlabel metal2 6692 11732 6692 11732 0 _037_
rlabel metal3 13552 11116 13552 11116 0 _038_
rlabel metal2 13300 13244 13300 13244 0 _039_
rlabel metal2 13692 12012 13692 12012 0 _040_
rlabel metal2 11228 13860 11228 13860 0 _041_
rlabel metal2 12180 13104 12180 13104 0 _042_
rlabel metal2 13132 13328 13132 13328 0 _043_
rlabel metal2 6804 8820 6804 8820 0 _044_
rlabel metal2 9212 8736 9212 8736 0 _045_
rlabel metal2 6860 8736 6860 8736 0 _046_
rlabel metal3 11816 13916 11816 13916 0 _047_
rlabel metal2 11900 12964 11900 12964 0 _048_
rlabel metal3 13188 13132 13188 13132 0 _049_
rlabel metal2 9044 13244 9044 13244 0 _050_
rlabel metal2 13244 7840 13244 7840 0 _051_
rlabel metal3 7672 8764 7672 8764 0 _052_
rlabel metal2 13692 10752 13692 10752 0 _053_
rlabel metal2 8876 10388 8876 10388 0 _054_
rlabel metal2 11844 8904 11844 8904 0 _055_
rlabel metal3 9576 10108 9576 10108 0 _056_
rlabel metal3 12740 9604 12740 9604 0 _057_
rlabel metal2 10332 11060 10332 11060 0 _058_
rlabel metal2 11228 9128 11228 9128 0 _059_
rlabel metal3 12572 10724 12572 10724 0 _060_
rlabel metal3 8624 10052 8624 10052 0 _061_
rlabel metal3 8288 10388 8288 10388 0 _062_
rlabel metal2 11788 9632 11788 9632 0 _063_
rlabel metal2 9212 8372 9212 8372 0 _064_
rlabel metal2 9884 9016 9884 9016 0 _065_
rlabel metal2 8400 10164 8400 10164 0 _066_
rlabel metal3 11228 8820 11228 8820 0 _067_
rlabel metal2 10500 11312 10500 11312 0 _068_
rlabel metal2 12348 10864 12348 10864 0 _069_
rlabel metal2 8820 12824 8820 12824 0 _070_
rlabel metal2 8848 8148 8848 8148 0 _071_
rlabel metal3 10388 10976 10388 10976 0 _072_
rlabel metal2 12124 9576 12124 9576 0 _073_
rlabel metal2 11396 11396 11396 11396 0 _074_
rlabel metal2 12768 11172 12768 11172 0 _075_
rlabel metal3 10808 9100 10808 9100 0 _076_
rlabel metal2 11452 8512 11452 8512 0 _077_
rlabel metal2 11480 12012 11480 12012 0 _078_
rlabel metal2 10108 12292 10108 12292 0 _079_
rlabel metal3 10346 11172 10346 11172 0 _080_
rlabel via2 10220 9044 10220 9044 0 _081_
rlabel metal2 11956 12880 11956 12880 0 _082_
rlabel metal3 8428 11676 8428 11676 0 _083_
rlabel metal3 12404 11228 12404 11228 0 _084_
rlabel metal2 10108 9716 10108 9716 0 _085_
rlabel metal3 7420 9996 7420 9996 0 _086_
rlabel metal2 10612 12964 10612 12964 0 _087_
rlabel metal2 13076 11984 13076 11984 0 _088_
rlabel metal2 6916 11788 6916 11788 0 _089_
rlabel metal3 7364 12460 7364 12460 0 _090_
rlabel metal2 6524 9996 6524 9996 0 _091_
rlabel metal3 11368 9212 11368 9212 0 _092_
rlabel metal2 12292 8764 12292 8764 0 _093_
rlabel metal2 12236 8680 12236 8680 0 _094_
rlabel metal2 12180 11396 12180 11396 0 _095_
rlabel metal2 11984 11452 11984 11452 0 _096_
rlabel metal3 1239 14140 1239 14140 0 clk
rlabel metal2 12628 10612 12628 10612 0 clknet_0_clk
rlabel metal2 11004 13160 11004 13160 0 clknet_1_0__leaf_clk
rlabel metal3 11816 14252 11816 14252 0 clknet_1_1__leaf_clk
rlabel metal2 12012 11032 12012 11032 0 dut47.count\[0\]
rlabel metal2 11564 10808 11564 10808 0 dut47.count\[1\]
rlabel metal2 8316 11312 8316 11312 0 dut47.count\[2\]
rlabel metal3 8512 9996 8512 9996 0 dut47.count\[3\]
rlabel metal2 5460 9184 5460 9184 0 net1
rlabel metal3 16240 8092 16240 8092 0 net10
rlabel metal2 12572 14672 12572 14672 0 net11
rlabel metal2 14084 14056 14084 14056 0 net12
rlabel metal2 10724 13496 10724 13496 0 net13
rlabel metal2 14196 11536 14196 11536 0 net14
rlabel metal3 16772 12292 16772 12292 0 net15
rlabel metal3 16576 8372 16576 8372 0 net16
rlabel metal2 7308 13496 7308 13496 0 net17
rlabel metal2 5572 12124 5572 12124 0 net18
rlabel metal3 10752 6804 10752 6804 0 net19
rlabel metal2 12404 14336 12404 14336 0 net2
rlabel metal2 13356 8316 13356 8316 0 net20
rlabel metal2 8820 2982 8820 2982 0 net21
rlabel metal3 5852 10444 5852 10444 0 net22
rlabel metal2 6356 8596 6356 8596 0 net23
rlabel metal2 13804 10556 13804 10556 0 net24
rlabel metal2 8708 18956 8708 18956 0 net25
rlabel metal3 623 18172 623 18172 0 net26
rlabel metal2 13664 13580 13664 13580 0 net3
rlabel metal2 9240 13244 9240 13244 0 net4
rlabel metal2 11900 3374 11900 3374 0 net5
rlabel metal2 7644 13580 7644 13580 0 net6
rlabel metal2 12292 2982 12292 2982 0 net7
rlabel metal2 5964 13104 5964 13104 0 net8
rlabel metal2 9856 2156 9856 2156 0 net9
rlabel metal3 679 9100 679 9100 0 segm[10]
rlabel metal2 12124 19873 12124 19873 0 segm[11]
rlabel metal2 13804 19677 13804 19677 0 segm[12]
rlabel metal2 9100 19873 9100 19873 0 segm[13]
rlabel metal2 11788 1491 11788 1491 0 segm[1]
rlabel metal3 679 13468 679 13468 0 segm[2]
rlabel metal2 11452 1099 11452 1099 0 segm[4]
rlabel metal3 679 12796 679 12796 0 segm[5]
rlabel metal2 9772 1211 9772 1211 0 segm[6]
rlabel metal3 20321 8092 20321 8092 0 segm[7]
rlabel metal2 12460 19677 12460 19677 0 segm[8]
rlabel metal2 13468 19873 13468 19873 0 segm[9]
rlabel metal2 10780 19873 10780 19873 0 sel[0]
rlabel metal3 20321 11452 20321 11452 0 sel[10]
rlabel metal2 20020 12628 20020 12628 0 sel[11]
rlabel metal2 20020 8820 20020 8820 0 sel[1]
rlabel metal3 707 13132 707 13132 0 sel[2]
rlabel metal3 679 11788 679 11788 0 sel[3]
rlabel metal2 11116 1015 11116 1015 0 sel[4]
rlabel metal2 20020 8400 20020 8400 0 sel[5]
rlabel metal2 8764 1099 8764 1099 0 sel[6]
rlabel metal3 679 10444 679 10444 0 sel[7]
rlabel metal3 679 8428 679 8428 0 sel[8]
rlabel metal2 20020 10556 20020 10556 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
