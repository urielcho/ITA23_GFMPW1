magic
tech gf180mcuD
magscale 1 10
timestamp 1699641367
<< metal1 >>
rect 18834 38558 18846 38610
rect 18898 38607 18910 38610
rect 19954 38607 19966 38610
rect 18898 38561 19966 38607
rect 18898 38558 18910 38561
rect 19954 38558 19966 38561
rect 20018 38558 20030 38610
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18062 38274 18114 38286
rect 18062 38210 18114 38222
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 17266 37998 17278 38050
rect 17330 37998 17342 38050
rect 21746 37998 21758 38050
rect 21810 37998 21822 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 19966 37938 20018 37950
rect 19966 37874 20018 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 20750 37490 20802 37502
rect 20750 37426 20802 37438
rect 19730 37214 19742 37266
rect 19794 37214 19806 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 40238 36370 40290 36382
rect 40238 36306 40290 36318
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 19506 27134 19518 27186
rect 19570 27134 19582 27186
rect 24322 27134 24334 27186
rect 24386 27134 24398 27186
rect 20414 27074 20466 27086
rect 24782 27074 24834 27086
rect 16706 27022 16718 27074
rect 16770 27022 16782 27074
rect 21522 27022 21534 27074
rect 21586 27022 21598 27074
rect 20414 27010 20466 27022
rect 24782 27010 24834 27022
rect 19854 26962 19906 26974
rect 17378 26910 17390 26962
rect 17442 26910 17454 26962
rect 22194 26910 22206 26962
rect 22258 26910 22270 26962
rect 19854 26898 19906 26910
rect 19742 26850 19794 26862
rect 19742 26786 19794 26798
rect 20078 26850 20130 26862
rect 20078 26786 20130 26798
rect 20750 26850 20802 26862
rect 20750 26786 20802 26798
rect 40238 26850 40290 26862
rect 40238 26786 40290 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 18062 26514 18114 26526
rect 18062 26450 18114 26462
rect 21982 26514 22034 26526
rect 21982 26450 22034 26462
rect 22206 26514 22258 26526
rect 22206 26450 22258 26462
rect 22990 26514 23042 26526
rect 22990 26450 23042 26462
rect 22318 26402 22370 26414
rect 19618 26350 19630 26402
rect 19682 26350 19694 26402
rect 22318 26338 22370 26350
rect 17950 26290 18002 26302
rect 13906 26238 13918 26290
rect 13970 26238 13982 26290
rect 17950 26226 18002 26238
rect 18286 26290 18338 26302
rect 18286 26226 18338 26238
rect 18510 26290 18562 26302
rect 22878 26290 22930 26302
rect 18946 26238 18958 26290
rect 19010 26238 19022 26290
rect 22642 26238 22654 26290
rect 22706 26238 22718 26290
rect 18510 26226 18562 26238
rect 22878 26226 22930 26238
rect 23102 26290 23154 26302
rect 23314 26238 23326 26290
rect 23378 26238 23390 26290
rect 37874 26238 37886 26290
rect 37938 26238 37950 26290
rect 23102 26226 23154 26238
rect 13134 26178 13186 26190
rect 17502 26178 17554 26190
rect 14578 26126 14590 26178
rect 14642 26126 14654 26178
rect 16706 26126 16718 26178
rect 16770 26126 16782 26178
rect 21746 26126 21758 26178
rect 21810 26126 21822 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 13134 26114 13186 26126
rect 17502 26114 17554 26126
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 1934 25618 1986 25630
rect 18510 25618 18562 25630
rect 40014 25618 40066 25630
rect 9986 25566 9998 25618
rect 10050 25566 10062 25618
rect 19394 25566 19406 25618
rect 19458 25566 19470 25618
rect 26898 25566 26910 25618
rect 26962 25566 26974 25618
rect 1934 25554 1986 25566
rect 18510 25554 18562 25566
rect 40014 25554 40066 25566
rect 13694 25506 13746 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 12898 25454 12910 25506
rect 12962 25454 12974 25506
rect 13694 25442 13746 25454
rect 13806 25506 13858 25518
rect 13806 25442 13858 25454
rect 15038 25506 15090 25518
rect 15038 25442 15090 25454
rect 15374 25506 15426 25518
rect 15374 25442 15426 25454
rect 16382 25506 16434 25518
rect 16382 25442 16434 25454
rect 16494 25506 16546 25518
rect 19854 25506 19906 25518
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 19282 25454 19294 25506
rect 19346 25454 19358 25506
rect 16494 25442 16546 25454
rect 19854 25442 19906 25454
rect 21198 25506 21250 25518
rect 23986 25454 23998 25506
rect 24050 25454 24062 25506
rect 27346 25454 27358 25506
rect 27410 25454 27422 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 21198 25442 21250 25454
rect 14030 25394 14082 25406
rect 12114 25342 12126 25394
rect 12178 25342 12190 25394
rect 14030 25330 14082 25342
rect 14142 25394 14194 25406
rect 14142 25330 14194 25342
rect 21422 25394 21474 25406
rect 21422 25330 21474 25342
rect 21534 25394 21586 25406
rect 24770 25342 24782 25394
rect 24834 25342 24846 25394
rect 21534 25330 21586 25342
rect 15262 25282 15314 25294
rect 15262 25218 15314 25230
rect 16270 25282 16322 25294
rect 16270 25218 16322 25230
rect 19518 25282 19570 25294
rect 19518 25218 19570 25230
rect 19742 25282 19794 25294
rect 28030 25282 28082 25294
rect 27570 25230 27582 25282
rect 27634 25230 27646 25282
rect 19742 25218 19794 25230
rect 28030 25218 28082 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 14030 24946 14082 24958
rect 14030 24882 14082 24894
rect 14254 24946 14306 24958
rect 14254 24882 14306 24894
rect 16046 24946 16098 24958
rect 16046 24882 16098 24894
rect 19854 24946 19906 24958
rect 19854 24882 19906 24894
rect 20190 24946 20242 24958
rect 20190 24882 20242 24894
rect 25566 24834 25618 24846
rect 21298 24782 21310 24834
rect 21362 24782 21374 24834
rect 25566 24770 25618 24782
rect 14366 24722 14418 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 13794 24670 13806 24722
rect 13858 24670 13870 24722
rect 14366 24658 14418 24670
rect 19742 24722 19794 24734
rect 19742 24658 19794 24670
rect 19966 24722 20018 24734
rect 19966 24658 20018 24670
rect 21646 24722 21698 24734
rect 21646 24658 21698 24670
rect 14814 24610 14866 24622
rect 10882 24558 10894 24610
rect 10946 24558 10958 24610
rect 13010 24558 13022 24610
rect 13074 24558 13086 24610
rect 14814 24546 14866 24558
rect 16158 24610 16210 24622
rect 16158 24546 16210 24558
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 25454 24498 25506 24510
rect 25454 24434 25506 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 19182 24162 19234 24174
rect 19182 24098 19234 24110
rect 1934 24050 1986 24062
rect 1934 23986 1986 23998
rect 12798 24050 12850 24062
rect 17054 24050 17106 24062
rect 24334 24050 24386 24062
rect 28366 24050 28418 24062
rect 13682 23998 13694 24050
rect 13746 23998 13758 24050
rect 21858 23998 21870 24050
rect 21922 23998 21934 24050
rect 27906 23998 27918 24050
rect 27970 23998 27982 24050
rect 12798 23986 12850 23998
rect 17054 23986 17106 23998
rect 24334 23986 24386 23998
rect 28366 23986 28418 23998
rect 18958 23938 19010 23950
rect 24110 23938 24162 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 16594 23886 16606 23938
rect 16658 23886 16670 23938
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 24658 23886 24670 23938
rect 24722 23886 24734 23938
rect 24994 23886 25006 23938
rect 25058 23886 25070 23938
rect 18958 23874 19010 23886
rect 24110 23874 24162 23886
rect 12686 23826 12738 23838
rect 12686 23762 12738 23774
rect 12910 23826 12962 23838
rect 20750 23826 20802 23838
rect 15810 23774 15822 23826
rect 15874 23774 15886 23826
rect 12910 23762 12962 23774
rect 20750 23762 20802 23774
rect 22094 23826 22146 23838
rect 25778 23774 25790 23826
rect 25842 23774 25854 23826
rect 22094 23762 22146 23774
rect 19294 23714 19346 23726
rect 19294 23650 19346 23662
rect 19518 23714 19570 23726
rect 19518 23650 19570 23662
rect 20414 23714 20466 23726
rect 20414 23650 20466 23662
rect 20638 23714 20690 23726
rect 23214 23714 23266 23726
rect 22418 23662 22430 23714
rect 22482 23662 22494 23714
rect 20638 23650 20690 23662
rect 23214 23650 23266 23662
rect 24222 23714 24274 23726
rect 24222 23650 24274 23662
rect 24446 23714 24498 23726
rect 24446 23650 24498 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 13918 23378 13970 23390
rect 25678 23378 25730 23390
rect 15810 23326 15822 23378
rect 15874 23326 15886 23378
rect 17378 23326 17390 23378
rect 17442 23326 17454 23378
rect 13918 23314 13970 23326
rect 25678 23314 25730 23326
rect 13806 23266 13858 23278
rect 13806 23202 13858 23214
rect 14142 23266 14194 23278
rect 14142 23202 14194 23214
rect 15486 23266 15538 23278
rect 23886 23266 23938 23278
rect 15698 23214 15710 23266
rect 15762 23214 15774 23266
rect 18274 23214 18286 23266
rect 18338 23214 18350 23266
rect 15486 23202 15538 23214
rect 23886 23202 23938 23214
rect 25454 23266 25506 23278
rect 25454 23202 25506 23214
rect 14366 23154 14418 23166
rect 18622 23154 18674 23166
rect 23102 23154 23154 23166
rect 25230 23154 25282 23166
rect 16258 23102 16270 23154
rect 16322 23102 16334 23154
rect 17602 23102 17614 23154
rect 17666 23102 17678 23154
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 23314 23102 23326 23154
rect 23378 23102 23390 23154
rect 14366 23090 14418 23102
rect 18622 23090 18674 23102
rect 23102 23090 23154 23102
rect 25230 23090 25282 23102
rect 25790 23154 25842 23166
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 25790 23090 25842 23102
rect 22430 23042 22482 23054
rect 19954 22990 19966 23042
rect 20018 22990 20030 23042
rect 22082 22990 22094 23042
rect 22146 22990 22158 23042
rect 22754 22990 22766 23042
rect 22818 22990 22830 23042
rect 22430 22978 22482 22990
rect 15934 22930 15986 22942
rect 15934 22866 15986 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 16270 22482 16322 22494
rect 16270 22418 16322 22430
rect 19070 22482 19122 22494
rect 25790 22482 25842 22494
rect 19394 22430 19406 22482
rect 19458 22430 19470 22482
rect 19070 22418 19122 22430
rect 25790 22418 25842 22430
rect 15934 22370 15986 22382
rect 15934 22306 15986 22318
rect 16046 22370 16098 22382
rect 16046 22306 16098 22318
rect 16494 22370 16546 22382
rect 16494 22306 16546 22318
rect 17166 22370 17218 22382
rect 17166 22306 17218 22318
rect 17278 22370 17330 22382
rect 17938 22318 17950 22370
rect 18002 22318 18014 22370
rect 19506 22318 19518 22370
rect 19570 22318 19582 22370
rect 20290 22318 20302 22370
rect 20354 22318 20366 22370
rect 23090 22318 23102 22370
rect 23154 22318 23166 22370
rect 23538 22318 23550 22370
rect 23602 22318 23614 22370
rect 26114 22318 26126 22370
rect 26178 22318 26190 22370
rect 17278 22306 17330 22318
rect 24558 22258 24610 22270
rect 18162 22206 18174 22258
rect 18226 22206 18238 22258
rect 18722 22206 18734 22258
rect 18786 22206 18798 22258
rect 19282 22206 19294 22258
rect 19346 22206 19358 22258
rect 21298 22206 21310 22258
rect 21362 22206 21374 22258
rect 24558 22194 24610 22206
rect 25678 22258 25730 22270
rect 25678 22194 25730 22206
rect 16830 22146 16882 22158
rect 25566 22146 25618 22158
rect 24994 22094 25006 22146
rect 25058 22094 25070 22146
rect 16830 22082 16882 22094
rect 25566 22082 25618 22094
rect 25902 22146 25954 22158
rect 25902 22082 25954 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 13470 21810 13522 21822
rect 13470 21746 13522 21758
rect 14142 21810 14194 21822
rect 14142 21746 14194 21758
rect 17950 21810 18002 21822
rect 25566 21810 25618 21822
rect 19058 21758 19070 21810
rect 19122 21758 19134 21810
rect 25218 21758 25230 21810
rect 25282 21758 25294 21810
rect 17950 21746 18002 21758
rect 25566 21746 25618 21758
rect 13246 21698 13298 21710
rect 13246 21634 13298 21646
rect 15150 21698 15202 21710
rect 15150 21634 15202 21646
rect 14926 21586 14978 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 12898 21534 12910 21586
rect 12962 21534 12974 21586
rect 13682 21534 13694 21586
rect 13746 21534 13758 21586
rect 14926 21522 14978 21534
rect 15262 21586 15314 21598
rect 18286 21586 18338 21598
rect 26014 21586 26066 21598
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 18834 21534 18846 21586
rect 18898 21534 18910 21586
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 15262 21522 15314 21534
rect 18286 21522 18338 21534
rect 26014 21522 26066 21534
rect 26238 21586 26290 21598
rect 26238 21522 26290 21534
rect 26574 21586 26626 21598
rect 26898 21534 26910 21586
rect 26962 21534 26974 21586
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 26574 21522 26626 21534
rect 17502 21474 17554 21486
rect 9986 21422 9998 21474
rect 10050 21422 10062 21474
rect 12114 21422 12126 21474
rect 12178 21422 12190 21474
rect 17502 21410 17554 21422
rect 18062 21474 18114 21486
rect 26462 21474 26514 21486
rect 30270 21474 30322 21486
rect 23314 21422 23326 21474
rect 23378 21422 23390 21474
rect 27682 21422 27694 21474
rect 27746 21422 27758 21474
rect 29810 21422 29822 21474
rect 29874 21422 29886 21474
rect 39890 21422 39902 21474
rect 39954 21422 39966 21474
rect 18062 21410 18114 21422
rect 26462 21410 26514 21422
rect 30270 21410 30322 21422
rect 1934 21362 1986 21374
rect 1934 21298 1986 21310
rect 13134 21362 13186 21374
rect 13134 21298 13186 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 15150 20914 15202 20926
rect 21982 20914 22034 20926
rect 40014 20914 40066 20926
rect 2034 20862 2046 20914
rect 2098 20862 2110 20914
rect 9986 20862 9998 20914
rect 10050 20862 10062 20914
rect 15698 20862 15710 20914
rect 15762 20862 15774 20914
rect 26898 20862 26910 20914
rect 26962 20862 26974 20914
rect 15150 20850 15202 20862
rect 21982 20850 22034 20862
rect 40014 20850 40066 20862
rect 13470 20802 13522 20814
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 12898 20750 12910 20802
rect 12962 20750 12974 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 22306 20750 22318 20802
rect 22370 20750 22382 20802
rect 22866 20750 22878 20802
rect 22930 20750 22942 20802
rect 23314 20750 23326 20802
rect 23378 20750 23390 20802
rect 29474 20750 29486 20802
rect 29538 20750 29550 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 13470 20738 13522 20750
rect 13806 20690 13858 20702
rect 12114 20638 12126 20690
rect 12178 20638 12190 20690
rect 13806 20626 13858 20638
rect 14030 20690 14082 20702
rect 29150 20690 29202 20702
rect 14354 20638 14366 20690
rect 14418 20638 14430 20690
rect 21522 20638 21534 20690
rect 21586 20638 21598 20690
rect 14030 20626 14082 20638
rect 29150 20626 29202 20638
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 14702 20578 14754 20590
rect 14702 20514 14754 20526
rect 29262 20578 29314 20590
rect 29262 20514 29314 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 12350 20242 12402 20254
rect 12350 20178 12402 20190
rect 18958 20242 19010 20254
rect 18958 20178 19010 20190
rect 19966 20242 20018 20254
rect 19966 20178 20018 20190
rect 23102 20242 23154 20254
rect 23102 20178 23154 20190
rect 12574 20130 12626 20142
rect 12574 20066 12626 20078
rect 12686 20130 12738 20142
rect 12686 20066 12738 20078
rect 19742 20130 19794 20142
rect 19742 20066 19794 20078
rect 20862 20130 20914 20142
rect 20862 20066 20914 20078
rect 24446 20130 24498 20142
rect 24446 20066 24498 20078
rect 24558 20130 24610 20142
rect 24558 20066 24610 20078
rect 24782 20130 24834 20142
rect 24782 20066 24834 20078
rect 25342 20130 25394 20142
rect 27346 20078 27358 20130
rect 27410 20078 27422 20130
rect 25342 20066 25394 20078
rect 18622 20018 18674 20030
rect 19518 20018 19570 20030
rect 22766 20018 22818 20030
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 15810 19966 15822 20018
rect 15874 19966 15886 20018
rect 16258 19966 16270 20018
rect 16322 19966 16334 20018
rect 19170 19966 19182 20018
rect 19234 19966 19246 20018
rect 20178 19966 20190 20018
rect 20242 19966 20254 20018
rect 21410 19966 21422 20018
rect 21474 19966 21486 20018
rect 22530 19966 22542 20018
rect 22594 19966 22606 20018
rect 18622 19954 18674 19966
rect 19518 19954 19570 19966
rect 22766 19954 22818 19966
rect 23774 20018 23826 20030
rect 23774 19954 23826 19966
rect 25118 20018 25170 20030
rect 25118 19954 25170 19966
rect 25454 20018 25506 20030
rect 25454 19954 25506 19966
rect 25790 20018 25842 20030
rect 26674 19966 26686 20018
rect 26738 19966 26750 20018
rect 25790 19954 25842 19966
rect 16606 19906 16658 19918
rect 23550 19906 23602 19918
rect 29934 19906 29986 19918
rect 13010 19854 13022 19906
rect 13074 19854 13086 19906
rect 15138 19854 15150 19906
rect 15202 19854 15214 19906
rect 18162 19854 18174 19906
rect 18226 19854 18238 19906
rect 21298 19854 21310 19906
rect 21362 19854 21374 19906
rect 29474 19854 29486 19906
rect 29538 19854 29550 19906
rect 16606 19842 16658 19854
rect 23550 19842 23602 19854
rect 29934 19842 29986 19854
rect 1934 19794 1986 19806
rect 1934 19730 1986 19742
rect 16270 19794 16322 19806
rect 16270 19730 16322 19742
rect 18846 19794 18898 19806
rect 18846 19730 18898 19742
rect 19630 19794 19682 19806
rect 19630 19730 19682 19742
rect 24110 19794 24162 19806
rect 24110 19730 24162 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 14926 19458 14978 19470
rect 14926 19394 14978 19406
rect 15262 19458 15314 19470
rect 15262 19394 15314 19406
rect 26350 19458 26402 19470
rect 26350 19394 26402 19406
rect 27022 19458 27074 19470
rect 27022 19394 27074 19406
rect 27134 19458 27186 19470
rect 27134 19394 27186 19406
rect 27358 19458 27410 19470
rect 27358 19394 27410 19406
rect 27470 19458 27522 19470
rect 27470 19394 27522 19406
rect 16158 19346 16210 19358
rect 24334 19346 24386 19358
rect 21858 19294 21870 19346
rect 21922 19294 21934 19346
rect 25106 19294 25118 19346
rect 25170 19294 25182 19346
rect 16158 19282 16210 19294
rect 24334 19282 24386 19294
rect 15038 19234 15090 19246
rect 20750 19234 20802 19246
rect 15474 19182 15486 19234
rect 15538 19182 15550 19234
rect 18050 19182 18062 19234
rect 18114 19182 18126 19234
rect 18498 19182 18510 19234
rect 18562 19182 18574 19234
rect 19170 19182 19182 19234
rect 19234 19182 19246 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 22530 19182 22542 19234
rect 22594 19182 22606 19234
rect 23762 19182 23774 19234
rect 23826 19182 23838 19234
rect 24098 19182 24110 19234
rect 24162 19182 24174 19234
rect 25778 19182 25790 19234
rect 25842 19182 25854 19234
rect 15038 19170 15090 19182
rect 20750 19170 20802 19182
rect 17726 19122 17778 19134
rect 26238 19122 26290 19134
rect 18722 19070 18734 19122
rect 18786 19070 18798 19122
rect 19730 19070 19742 19122
rect 19794 19070 19806 19122
rect 20402 19070 20414 19122
rect 20466 19070 20478 19122
rect 21634 19070 21646 19122
rect 21698 19070 21710 19122
rect 17726 19058 17778 19070
rect 26238 19058 26290 19070
rect 17278 19010 17330 19022
rect 16930 18958 16942 19010
rect 16994 18958 17006 19010
rect 17278 18946 17330 18958
rect 17838 19010 17890 19022
rect 20078 19010 20130 19022
rect 19394 18958 19406 19010
rect 19458 18958 19470 19010
rect 17838 18946 17890 18958
rect 20078 18946 20130 18958
rect 24670 19010 24722 19022
rect 24670 18946 24722 18958
rect 26014 19010 26066 19022
rect 26014 18946 26066 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 20750 18674 20802 18686
rect 17714 18622 17726 18674
rect 17778 18622 17790 18674
rect 20750 18610 20802 18622
rect 21310 18674 21362 18686
rect 21310 18610 21362 18622
rect 21198 18562 21250 18574
rect 21970 18510 21982 18562
rect 22034 18510 22046 18562
rect 23874 18510 23886 18562
rect 23938 18510 23950 18562
rect 21198 18498 21250 18510
rect 16382 18450 16434 18462
rect 19070 18450 19122 18462
rect 21534 18450 21586 18462
rect 24334 18450 24386 18462
rect 28030 18450 28082 18462
rect 16034 18398 16046 18450
rect 16098 18398 16110 18450
rect 17490 18398 17502 18450
rect 17554 18398 17566 18450
rect 18610 18398 18622 18450
rect 18674 18398 18686 18450
rect 19282 18398 19294 18450
rect 19346 18398 19358 18450
rect 22306 18398 22318 18450
rect 22370 18398 22382 18450
rect 22754 18398 22766 18450
rect 22818 18398 22830 18450
rect 23314 18398 23326 18450
rect 23378 18398 23390 18450
rect 27682 18398 27694 18450
rect 27746 18398 27758 18450
rect 16382 18386 16434 18398
rect 19070 18386 19122 18398
rect 21534 18386 21586 18398
rect 24334 18386 24386 18398
rect 28030 18386 28082 18398
rect 28478 18450 28530 18462
rect 28690 18398 28702 18450
rect 28754 18398 28766 18450
rect 37874 18398 37886 18450
rect 37938 18398 37950 18450
rect 28478 18386 28530 18398
rect 19854 18338 19906 18350
rect 18274 18286 18286 18338
rect 18338 18286 18350 18338
rect 19854 18274 19906 18286
rect 20190 18338 20242 18350
rect 23650 18286 23662 18338
rect 23714 18286 23726 18338
rect 20190 18274 20242 18286
rect 16046 18226 16098 18238
rect 16046 18162 16098 18174
rect 27694 18226 27746 18238
rect 27694 18162 27746 18174
rect 28366 18226 28418 18238
rect 28366 18162 28418 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 18062 17890 18114 17902
rect 18062 17826 18114 17838
rect 18846 17890 18898 17902
rect 18846 17826 18898 17838
rect 20638 17890 20690 17902
rect 20638 17826 20690 17838
rect 1934 17778 1986 17790
rect 1934 17714 1986 17726
rect 14478 17778 14530 17790
rect 14478 17714 14530 17726
rect 17054 17778 17106 17790
rect 40014 17778 40066 17790
rect 23762 17726 23774 17778
rect 23826 17726 23838 17778
rect 17054 17714 17106 17726
rect 40014 17714 40066 17726
rect 12574 17666 12626 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 12574 17602 12626 17614
rect 12910 17666 12962 17678
rect 12910 17602 12962 17614
rect 13358 17666 13410 17678
rect 13358 17602 13410 17614
rect 13806 17666 13858 17678
rect 13806 17602 13858 17614
rect 13918 17666 13970 17678
rect 26014 17666 26066 17678
rect 18050 17614 18062 17666
rect 18114 17614 18126 17666
rect 22978 17614 22990 17666
rect 23042 17614 23054 17666
rect 24098 17614 24110 17666
rect 24162 17614 24174 17666
rect 24434 17614 24446 17666
rect 24498 17614 24510 17666
rect 13918 17602 13970 17614
rect 26014 17602 26066 17614
rect 26462 17666 26514 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 26462 17602 26514 17614
rect 12798 17554 12850 17566
rect 12798 17490 12850 17502
rect 17390 17554 17442 17566
rect 18398 17554 18450 17566
rect 17714 17502 17726 17554
rect 17778 17502 17790 17554
rect 17390 17490 17442 17502
rect 18398 17490 18450 17502
rect 18734 17554 18786 17566
rect 18734 17490 18786 17502
rect 20750 17554 20802 17566
rect 22194 17502 22206 17554
rect 22258 17502 22270 17554
rect 23202 17502 23214 17554
rect 23266 17502 23278 17554
rect 20750 17490 20802 17502
rect 13582 17442 13634 17454
rect 13582 17378 13634 17390
rect 22542 17442 22594 17454
rect 26574 17442 26626 17454
rect 24770 17390 24782 17442
rect 24834 17390 24846 17442
rect 22542 17378 22594 17390
rect 26574 17378 26626 17390
rect 26686 17442 26738 17454
rect 26686 17378 26738 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 18846 17106 18898 17118
rect 18846 17042 18898 17054
rect 25566 17106 25618 17118
rect 25566 17042 25618 17054
rect 18174 16994 18226 17006
rect 19854 16994 19906 17006
rect 12450 16942 12462 16994
rect 12514 16942 12526 16994
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 18498 16942 18510 16994
rect 18562 16942 18574 16994
rect 18174 16930 18226 16942
rect 19854 16930 19906 16942
rect 19966 16994 20018 17006
rect 19966 16930 20018 16942
rect 21086 16994 21138 17006
rect 21086 16930 21138 16942
rect 21310 16994 21362 17006
rect 21310 16930 21362 16942
rect 25790 16994 25842 17006
rect 27682 16942 27694 16994
rect 27746 16942 27758 16994
rect 25790 16930 25842 16942
rect 17950 16882 18002 16894
rect 20190 16882 20242 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 13234 16830 13246 16882
rect 13298 16830 13310 16882
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 19170 16830 19182 16882
rect 19234 16830 19246 16882
rect 17950 16818 18002 16830
rect 20190 16818 20242 16830
rect 20638 16882 20690 16894
rect 30270 16882 30322 16894
rect 23762 16830 23774 16882
rect 23826 16830 23838 16882
rect 27010 16830 27022 16882
rect 27074 16830 27086 16882
rect 20638 16818 20690 16830
rect 30270 16818 30322 16830
rect 19518 16770 19570 16782
rect 10322 16718 10334 16770
rect 10386 16718 10398 16770
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 19518 16706 19570 16718
rect 20862 16770 20914 16782
rect 20862 16706 20914 16718
rect 23438 16770 23490 16782
rect 25678 16770 25730 16782
rect 23650 16718 23662 16770
rect 23714 16718 23726 16770
rect 29810 16718 29822 16770
rect 29874 16718 29886 16770
rect 23438 16706 23490 16718
rect 25678 16706 25730 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 17614 16658 17666 16670
rect 17614 16594 17666 16606
rect 19182 16658 19234 16670
rect 19182 16594 19234 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 25790 16210 25842 16222
rect 9986 16158 9998 16210
rect 10050 16158 10062 16210
rect 23650 16158 23662 16210
rect 23714 16158 23726 16210
rect 25790 16146 25842 16158
rect 13806 16098 13858 16110
rect 12898 16046 12910 16098
rect 12962 16046 12974 16098
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 13806 16034 13858 16046
rect 14030 16098 14082 16110
rect 16382 16098 16434 16110
rect 14690 16046 14702 16098
rect 14754 16046 14766 16098
rect 16818 16046 16830 16098
rect 16882 16046 16894 16098
rect 17154 16046 17166 16098
rect 17218 16046 17230 16098
rect 22978 16046 22990 16098
rect 23042 16046 23054 16098
rect 26562 16046 26574 16098
rect 26626 16046 26638 16098
rect 14030 16034 14082 16046
rect 16382 16034 16434 16046
rect 14366 15986 14418 15998
rect 12114 15934 12126 15986
rect 12178 15934 12190 15986
rect 14366 15922 14418 15934
rect 14478 15986 14530 15998
rect 14478 15922 14530 15934
rect 13918 15874 13970 15886
rect 13918 15810 13970 15822
rect 16494 15874 16546 15886
rect 16494 15810 16546 15822
rect 16606 15874 16658 15886
rect 27134 15874 27186 15886
rect 26338 15822 26350 15874
rect 26402 15822 26414 15874
rect 16606 15810 16658 15822
rect 27134 15810 27186 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 13134 15538 13186 15550
rect 13134 15474 13186 15486
rect 17502 15538 17554 15550
rect 17502 15474 17554 15486
rect 20738 15374 20750 15426
rect 20802 15374 20814 15426
rect 26002 15374 26014 15426
rect 26066 15374 26078 15426
rect 23326 15314 23378 15326
rect 28590 15314 28642 15326
rect 13906 15262 13918 15314
rect 13970 15262 13982 15314
rect 20066 15262 20078 15314
rect 20130 15262 20142 15314
rect 25330 15262 25342 15314
rect 25394 15262 25406 15314
rect 23326 15250 23378 15262
rect 28590 15250 28642 15262
rect 14690 15150 14702 15202
rect 14754 15150 14766 15202
rect 16818 15150 16830 15202
rect 16882 15150 16894 15202
rect 22866 15150 22878 15202
rect 22930 15150 22942 15202
rect 28130 15150 28142 15202
rect 28194 15150 28206 15202
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 15710 14754 15762 14766
rect 15710 14690 15762 14702
rect 15822 14642 15874 14654
rect 18610 14590 18622 14642
rect 18674 14590 18686 14642
rect 20738 14590 20750 14642
rect 20802 14590 20814 14642
rect 15822 14578 15874 14590
rect 17614 14530 17666 14542
rect 17826 14478 17838 14530
rect 17890 14478 17902 14530
rect 17614 14466 17666 14478
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 26798 4114 26850 4126
rect 26798 4050 26850 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 24782 3666 24834 3678
rect 24782 3602 24834 3614
rect 17042 3502 17054 3554
rect 17106 3502 17118 3554
rect 27122 3502 27134 3554
rect 27186 3502 27198 3554
rect 18062 3330 18114 3342
rect 18062 3266 18114 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 18846 38558 18898 38610
rect 19966 38558 20018 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18062 38222 18114 38274
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 17278 37998 17330 38050
rect 21758 37998 21810 38050
rect 24558 37998 24610 38050
rect 19966 37886 20018 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 20750 37438 20802 37490
rect 19742 37214 19794 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 1710 36318 1762 36370
rect 40238 36318 40290 36370
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 19518 27134 19570 27186
rect 24334 27134 24386 27186
rect 16718 27022 16770 27074
rect 20414 27022 20466 27074
rect 21534 27022 21586 27074
rect 24782 27022 24834 27074
rect 17390 26910 17442 26962
rect 19854 26910 19906 26962
rect 22206 26910 22258 26962
rect 19742 26798 19794 26850
rect 20078 26798 20130 26850
rect 20750 26798 20802 26850
rect 40238 26798 40290 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 18062 26462 18114 26514
rect 21982 26462 22034 26514
rect 22206 26462 22258 26514
rect 22990 26462 23042 26514
rect 19630 26350 19682 26402
rect 22318 26350 22370 26402
rect 13918 26238 13970 26290
rect 17950 26238 18002 26290
rect 18286 26238 18338 26290
rect 18510 26238 18562 26290
rect 18958 26238 19010 26290
rect 22654 26238 22706 26290
rect 22878 26238 22930 26290
rect 23102 26238 23154 26290
rect 23326 26238 23378 26290
rect 37886 26238 37938 26290
rect 13134 26126 13186 26178
rect 14590 26126 14642 26178
rect 16718 26126 16770 26178
rect 17502 26126 17554 26178
rect 21758 26126 21810 26178
rect 39902 26126 39954 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 1934 25566 1986 25618
rect 9998 25566 10050 25618
rect 18510 25566 18562 25618
rect 19406 25566 19458 25618
rect 26910 25566 26962 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 12910 25454 12962 25506
rect 13694 25454 13746 25506
rect 13806 25454 13858 25506
rect 15038 25454 15090 25506
rect 15374 25454 15426 25506
rect 16382 25454 16434 25506
rect 16494 25454 16546 25506
rect 16830 25454 16882 25506
rect 19294 25454 19346 25506
rect 19854 25454 19906 25506
rect 21198 25454 21250 25506
rect 23998 25454 24050 25506
rect 27358 25454 27410 25506
rect 37662 25454 37714 25506
rect 12126 25342 12178 25394
rect 14030 25342 14082 25394
rect 14142 25342 14194 25394
rect 21422 25342 21474 25394
rect 21534 25342 21586 25394
rect 24782 25342 24834 25394
rect 15262 25230 15314 25282
rect 16270 25230 16322 25282
rect 19518 25230 19570 25282
rect 19742 25230 19794 25282
rect 27582 25230 27634 25282
rect 28030 25230 28082 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 14030 24894 14082 24946
rect 14254 24894 14306 24946
rect 16046 24894 16098 24946
rect 19854 24894 19906 24946
rect 20190 24894 20242 24946
rect 21310 24782 21362 24834
rect 25566 24782 25618 24834
rect 4286 24670 4338 24722
rect 13806 24670 13858 24722
rect 14366 24670 14418 24722
rect 19742 24670 19794 24722
rect 19966 24670 20018 24722
rect 21646 24670 21698 24722
rect 10894 24558 10946 24610
rect 13022 24558 13074 24610
rect 14814 24558 14866 24610
rect 16158 24558 16210 24610
rect 1934 24446 1986 24498
rect 25454 24446 25506 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 19182 24110 19234 24162
rect 1934 23998 1986 24050
rect 12798 23998 12850 24050
rect 13694 23998 13746 24050
rect 17054 23998 17106 24050
rect 21870 23998 21922 24050
rect 24334 23998 24386 24050
rect 27918 23998 27970 24050
rect 28366 23998 28418 24050
rect 4286 23886 4338 23938
rect 16606 23886 16658 23938
rect 18958 23886 19010 23938
rect 22654 23886 22706 23938
rect 24110 23886 24162 23938
rect 24670 23886 24722 23938
rect 25006 23886 25058 23938
rect 12686 23774 12738 23826
rect 12910 23774 12962 23826
rect 15822 23774 15874 23826
rect 20750 23774 20802 23826
rect 22094 23774 22146 23826
rect 25790 23774 25842 23826
rect 19294 23662 19346 23714
rect 19518 23662 19570 23714
rect 20414 23662 20466 23714
rect 20638 23662 20690 23714
rect 22430 23662 22482 23714
rect 23214 23662 23266 23714
rect 24222 23662 24274 23714
rect 24446 23662 24498 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 13918 23326 13970 23378
rect 15822 23326 15874 23378
rect 17390 23326 17442 23378
rect 25678 23326 25730 23378
rect 13806 23214 13858 23266
rect 14142 23214 14194 23266
rect 15486 23214 15538 23266
rect 15710 23214 15762 23266
rect 18286 23214 18338 23266
rect 23886 23214 23938 23266
rect 25454 23214 25506 23266
rect 14366 23102 14418 23154
rect 16270 23102 16322 23154
rect 17614 23102 17666 23154
rect 18622 23102 18674 23154
rect 19182 23102 19234 23154
rect 23102 23102 23154 23154
rect 23326 23102 23378 23154
rect 25230 23102 25282 23154
rect 25790 23102 25842 23154
rect 37662 23102 37714 23154
rect 19966 22990 20018 23042
rect 22094 22990 22146 23042
rect 22430 22990 22482 23042
rect 22766 22990 22818 23042
rect 15934 22878 15986 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16270 22430 16322 22482
rect 19070 22430 19122 22482
rect 19406 22430 19458 22482
rect 25790 22430 25842 22482
rect 15934 22318 15986 22370
rect 16046 22318 16098 22370
rect 16494 22318 16546 22370
rect 17166 22318 17218 22370
rect 17278 22318 17330 22370
rect 17950 22318 18002 22370
rect 19518 22318 19570 22370
rect 20302 22318 20354 22370
rect 23102 22318 23154 22370
rect 23550 22318 23602 22370
rect 26126 22318 26178 22370
rect 18174 22206 18226 22258
rect 18734 22206 18786 22258
rect 19294 22206 19346 22258
rect 21310 22206 21362 22258
rect 24558 22206 24610 22258
rect 25678 22206 25730 22258
rect 16830 22094 16882 22146
rect 25006 22094 25058 22146
rect 25566 22094 25618 22146
rect 25902 22094 25954 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13470 21758 13522 21810
rect 14142 21758 14194 21810
rect 17950 21758 18002 21810
rect 19070 21758 19122 21810
rect 25230 21758 25282 21810
rect 25566 21758 25618 21810
rect 13246 21646 13298 21698
rect 15150 21646 15202 21698
rect 4286 21534 4338 21586
rect 12910 21534 12962 21586
rect 13694 21534 13746 21586
rect 14926 21534 14978 21586
rect 15262 21534 15314 21586
rect 17838 21534 17890 21586
rect 18286 21534 18338 21586
rect 18846 21534 18898 21586
rect 19406 21534 19458 21586
rect 26014 21534 26066 21586
rect 26238 21534 26290 21586
rect 26574 21534 26626 21586
rect 26910 21534 26962 21586
rect 37886 21534 37938 21586
rect 9998 21422 10050 21474
rect 12126 21422 12178 21474
rect 17502 21422 17554 21474
rect 18062 21422 18114 21474
rect 23326 21422 23378 21474
rect 26462 21422 26514 21474
rect 27694 21422 27746 21474
rect 29822 21422 29874 21474
rect 30270 21422 30322 21474
rect 39902 21422 39954 21474
rect 1934 21310 1986 21362
rect 13134 21310 13186 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 2046 20862 2098 20914
rect 9998 20862 10050 20914
rect 15150 20862 15202 20914
rect 15710 20862 15762 20914
rect 21982 20862 22034 20914
rect 26910 20862 26962 20914
rect 40014 20862 40066 20914
rect 4286 20750 4338 20802
rect 12910 20750 12962 20802
rect 13470 20750 13522 20802
rect 20078 20750 20130 20802
rect 21310 20750 21362 20802
rect 22318 20750 22370 20802
rect 22878 20750 22930 20802
rect 23326 20750 23378 20802
rect 29486 20750 29538 20802
rect 37662 20750 37714 20802
rect 12126 20638 12178 20690
rect 13806 20638 13858 20690
rect 14030 20638 14082 20690
rect 14366 20638 14418 20690
rect 21534 20638 21586 20690
rect 29150 20638 29202 20690
rect 13582 20526 13634 20578
rect 14702 20526 14754 20578
rect 29262 20526 29314 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 12350 20190 12402 20242
rect 18958 20190 19010 20242
rect 19966 20190 20018 20242
rect 23102 20190 23154 20242
rect 12574 20078 12626 20130
rect 12686 20078 12738 20130
rect 19742 20078 19794 20130
rect 20862 20078 20914 20130
rect 24446 20078 24498 20130
rect 24558 20078 24610 20130
rect 24782 20078 24834 20130
rect 25342 20078 25394 20130
rect 27358 20078 27410 20130
rect 4286 19966 4338 20018
rect 15822 19966 15874 20018
rect 16270 19966 16322 20018
rect 18622 19966 18674 20018
rect 19182 19966 19234 20018
rect 19518 19966 19570 20018
rect 20190 19966 20242 20018
rect 21422 19966 21474 20018
rect 22542 19966 22594 20018
rect 22766 19966 22818 20018
rect 23774 19966 23826 20018
rect 25118 19966 25170 20018
rect 25454 19966 25506 20018
rect 25790 19966 25842 20018
rect 26686 19966 26738 20018
rect 13022 19854 13074 19906
rect 15150 19854 15202 19906
rect 16606 19854 16658 19906
rect 18174 19854 18226 19906
rect 21310 19854 21362 19906
rect 23550 19854 23602 19906
rect 29486 19854 29538 19906
rect 29934 19854 29986 19906
rect 1934 19742 1986 19794
rect 16270 19742 16322 19794
rect 18846 19742 18898 19794
rect 19630 19742 19682 19794
rect 24110 19742 24162 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 14926 19406 14978 19458
rect 15262 19406 15314 19458
rect 26350 19406 26402 19458
rect 27022 19406 27074 19458
rect 27134 19406 27186 19458
rect 27358 19406 27410 19458
rect 27470 19406 27522 19458
rect 16158 19294 16210 19346
rect 21870 19294 21922 19346
rect 24334 19294 24386 19346
rect 25118 19294 25170 19346
rect 15038 19182 15090 19234
rect 15486 19182 15538 19234
rect 18062 19182 18114 19234
rect 18510 19182 18562 19234
rect 19182 19182 19234 19234
rect 20750 19182 20802 19234
rect 21534 19182 21586 19234
rect 22542 19182 22594 19234
rect 23774 19182 23826 19234
rect 24110 19182 24162 19234
rect 25790 19182 25842 19234
rect 17726 19070 17778 19122
rect 18734 19070 18786 19122
rect 19742 19070 19794 19122
rect 20414 19070 20466 19122
rect 21646 19070 21698 19122
rect 26238 19070 26290 19122
rect 16942 18958 16994 19010
rect 17278 18958 17330 19010
rect 17838 18958 17890 19010
rect 19406 18958 19458 19010
rect 20078 18958 20130 19010
rect 24670 18958 24722 19010
rect 26014 18958 26066 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 17726 18622 17778 18674
rect 20750 18622 20802 18674
rect 21310 18622 21362 18674
rect 21198 18510 21250 18562
rect 21982 18510 22034 18562
rect 23886 18510 23938 18562
rect 16046 18398 16098 18450
rect 16382 18398 16434 18450
rect 17502 18398 17554 18450
rect 18622 18398 18674 18450
rect 19070 18398 19122 18450
rect 19294 18398 19346 18450
rect 21534 18398 21586 18450
rect 22318 18398 22370 18450
rect 22766 18398 22818 18450
rect 23326 18398 23378 18450
rect 24334 18398 24386 18450
rect 27694 18398 27746 18450
rect 28030 18398 28082 18450
rect 28478 18398 28530 18450
rect 28702 18398 28754 18450
rect 37886 18398 37938 18450
rect 18286 18286 18338 18338
rect 19854 18286 19906 18338
rect 20190 18286 20242 18338
rect 23662 18286 23714 18338
rect 16046 18174 16098 18226
rect 27694 18174 27746 18226
rect 28366 18174 28418 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 18062 17838 18114 17890
rect 18846 17838 18898 17890
rect 20638 17838 20690 17890
rect 1934 17726 1986 17778
rect 14478 17726 14530 17778
rect 17054 17726 17106 17778
rect 23774 17726 23826 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 12574 17614 12626 17666
rect 12910 17614 12962 17666
rect 13358 17614 13410 17666
rect 13806 17614 13858 17666
rect 13918 17614 13970 17666
rect 18062 17614 18114 17666
rect 22990 17614 23042 17666
rect 24110 17614 24162 17666
rect 24446 17614 24498 17666
rect 26014 17614 26066 17666
rect 26462 17614 26514 17666
rect 37662 17614 37714 17666
rect 12798 17502 12850 17554
rect 17390 17502 17442 17554
rect 17726 17502 17778 17554
rect 18398 17502 18450 17554
rect 18734 17502 18786 17554
rect 20750 17502 20802 17554
rect 22206 17502 22258 17554
rect 23214 17502 23266 17554
rect 13582 17390 13634 17442
rect 22542 17390 22594 17442
rect 24782 17390 24834 17442
rect 26574 17390 26626 17442
rect 26686 17390 26738 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 18846 17054 18898 17106
rect 25566 17054 25618 17106
rect 12462 16942 12514 16994
rect 14702 16942 14754 16994
rect 18174 16942 18226 16994
rect 18510 16942 18562 16994
rect 19854 16942 19906 16994
rect 19966 16942 20018 16994
rect 21086 16942 21138 16994
rect 21310 16942 21362 16994
rect 25790 16942 25842 16994
rect 27694 16942 27746 16994
rect 4286 16830 4338 16882
rect 13246 16830 13298 16882
rect 14030 16830 14082 16882
rect 17950 16830 18002 16882
rect 19182 16830 19234 16882
rect 20190 16830 20242 16882
rect 20638 16830 20690 16882
rect 23774 16830 23826 16882
rect 27022 16830 27074 16882
rect 30270 16830 30322 16882
rect 10334 16718 10386 16770
rect 16830 16718 16882 16770
rect 19518 16718 19570 16770
rect 20862 16718 20914 16770
rect 23438 16718 23490 16770
rect 23662 16718 23714 16770
rect 25678 16718 25730 16770
rect 29822 16718 29874 16770
rect 1934 16606 1986 16658
rect 17614 16606 17666 16658
rect 19182 16606 19234 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 9998 16158 10050 16210
rect 23662 16158 23714 16210
rect 25790 16158 25842 16210
rect 12910 16046 12962 16098
rect 13470 16046 13522 16098
rect 13806 16046 13858 16098
rect 14030 16046 14082 16098
rect 14702 16046 14754 16098
rect 16382 16046 16434 16098
rect 16830 16046 16882 16098
rect 17166 16046 17218 16098
rect 22990 16046 23042 16098
rect 26574 16046 26626 16098
rect 12126 15934 12178 15986
rect 14366 15934 14418 15986
rect 14478 15934 14530 15986
rect 13918 15822 13970 15874
rect 16494 15822 16546 15874
rect 16606 15822 16658 15874
rect 26350 15822 26402 15874
rect 27134 15822 27186 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 13134 15486 13186 15538
rect 17502 15486 17554 15538
rect 20750 15374 20802 15426
rect 26014 15374 26066 15426
rect 13918 15262 13970 15314
rect 20078 15262 20130 15314
rect 23326 15262 23378 15314
rect 25342 15262 25394 15314
rect 28590 15262 28642 15314
rect 14702 15150 14754 15202
rect 16830 15150 16882 15202
rect 22878 15150 22930 15202
rect 28142 15150 28194 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 15710 14702 15762 14754
rect 15822 14590 15874 14642
rect 18622 14590 18674 14642
rect 20750 14590 20802 14642
rect 17614 14478 17666 14530
rect 17838 14478 17890 14530
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 25790 4286 25842 4338
rect 26798 4062 26850 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 24782 3614 24834 3666
rect 17054 3502 17106 3554
rect 27134 3502 27186 3554
rect 18062 3278 18114 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16800 41200 16912 42000
rect 18816 41200 18928 42000
rect 19488 41200 19600 42000
rect 21504 41200 21616 42000
rect 24192 41200 24304 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 16828 38276 16884 41200
rect 18844 38610 18900 41200
rect 18844 38558 18846 38610
rect 18898 38558 18900 38610
rect 18844 38546 18900 38558
rect 16828 38210 16884 38220
rect 18060 38276 18116 38286
rect 18060 38182 18116 38220
rect 17276 38050 17332 38062
rect 17276 37998 17278 38050
rect 17330 37998 17332 38050
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1708 36372 1764 36382
rect 1708 36278 1764 36316
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 16716 27074 16772 27086
rect 16716 27022 16718 27074
rect 16770 27022 16772 27074
rect 4172 26964 4228 26974
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 4172 21476 4228 26908
rect 16716 26908 16772 27022
rect 16716 26852 16996 26908
rect 13916 26290 13972 26302
rect 13916 26238 13918 26290
rect 13970 26238 13972 26290
rect 13132 26180 13188 26190
rect 12908 26124 13132 26180
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 9996 25620 10052 25630
rect 9996 25526 10052 25564
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 12908 25506 12964 26124
rect 13132 26086 13188 26124
rect 13916 26180 13972 26238
rect 16716 26292 16772 26302
rect 13804 25732 13860 25742
rect 12908 25454 12910 25506
rect 12962 25454 12964 25506
rect 12908 25442 12964 25454
rect 13692 25506 13748 25518
rect 13692 25454 13694 25506
rect 13746 25454 13748 25506
rect 12124 25396 12180 25406
rect 12124 25302 12180 25340
rect 12684 25284 12740 25294
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 10892 24612 10948 24622
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 10892 24164 10948 24556
rect 10892 24098 10948 24108
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 12684 23826 12740 25228
rect 13692 25284 13748 25454
rect 13804 25506 13860 25676
rect 13804 25454 13806 25506
rect 13858 25454 13860 25506
rect 13804 25442 13860 25454
rect 13692 25218 13748 25228
rect 13804 24724 13860 24734
rect 13916 24724 13972 26124
rect 14588 26180 14644 26190
rect 16716 26180 16772 26236
rect 14588 26178 15092 26180
rect 14588 26126 14590 26178
rect 14642 26126 15092 26178
rect 14588 26124 15092 26126
rect 14588 26114 14644 26124
rect 14252 25620 14308 25630
rect 14028 25396 14084 25406
rect 14028 25302 14084 25340
rect 14140 25394 14196 25406
rect 14140 25342 14142 25394
rect 14194 25342 14196 25394
rect 14028 24948 14084 24958
rect 14140 24948 14196 25342
rect 14028 24946 14196 24948
rect 14028 24894 14030 24946
rect 14082 24894 14196 24946
rect 14028 24892 14196 24894
rect 14252 24946 14308 25564
rect 15036 25506 15092 26124
rect 16492 26178 16772 26180
rect 16492 26126 16718 26178
rect 16770 26126 16772 26178
rect 16492 26124 16772 26126
rect 15036 25454 15038 25506
rect 15090 25454 15092 25506
rect 15036 25442 15092 25454
rect 15372 25508 15428 25518
rect 16380 25508 16436 25518
rect 15372 25506 16436 25508
rect 15372 25454 15374 25506
rect 15426 25454 16382 25506
rect 16434 25454 16436 25506
rect 15372 25452 16436 25454
rect 15372 25442 15428 25452
rect 16380 25442 16436 25452
rect 16492 25506 16548 26124
rect 16716 26114 16772 26124
rect 16940 26180 16996 26852
rect 17276 26292 17332 37998
rect 19516 37492 19572 41200
rect 19964 38610 20020 38622
rect 19964 38558 19966 38610
rect 20018 38558 20020 38610
rect 19964 37938 20020 38558
rect 21532 38276 21588 41200
rect 21532 38210 21588 38220
rect 22428 38276 22484 38286
rect 22428 38182 22484 38220
rect 24220 38276 24276 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 24220 38210 24276 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 19964 37886 19966 37938
rect 20018 37886 20020 37938
rect 19964 37874 20020 37886
rect 21756 38050 21812 38062
rect 21756 37998 21758 38050
rect 21810 37998 21812 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19516 37426 19572 37436
rect 20748 37492 20804 37502
rect 20748 37398 20804 37436
rect 19740 37268 19796 37278
rect 19516 37266 19796 37268
rect 19516 37214 19742 37266
rect 19794 37214 19796 37266
rect 19516 37212 19796 37214
rect 19516 27186 19572 37212
rect 19740 37202 19796 37212
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 27134 19518 27186
rect 19570 27134 19572 27186
rect 17388 26964 17444 26974
rect 17388 26962 18116 26964
rect 17388 26910 17390 26962
rect 17442 26910 18116 26962
rect 17388 26908 18116 26910
rect 17388 26898 17444 26908
rect 18060 26514 18116 26908
rect 18060 26462 18062 26514
rect 18114 26462 18116 26514
rect 18060 26450 18116 26462
rect 18956 26852 19012 26862
rect 17276 26226 17332 26236
rect 17948 26290 18004 26302
rect 17948 26238 17950 26290
rect 18002 26238 18004 26290
rect 16492 25454 16494 25506
rect 16546 25454 16548 25506
rect 16492 25442 16548 25454
rect 16828 25506 16884 25518
rect 16828 25454 16830 25506
rect 16882 25454 16884 25506
rect 14252 24894 14254 24946
rect 14306 24894 14308 24946
rect 14028 24882 14084 24892
rect 14252 24882 14308 24894
rect 15148 25284 15204 25294
rect 14364 24724 14420 24734
rect 13804 24722 13972 24724
rect 13804 24670 13806 24722
rect 13858 24670 13972 24722
rect 13804 24668 13972 24670
rect 13804 24658 13860 24668
rect 13020 24612 13076 24622
rect 12796 24610 13076 24612
rect 12796 24558 13022 24610
rect 13074 24558 13076 24610
rect 12796 24556 13076 24558
rect 12796 24050 12852 24556
rect 13020 24546 13076 24556
rect 13916 24612 13972 24668
rect 13916 24546 13972 24556
rect 14140 24722 14420 24724
rect 14140 24670 14366 24722
rect 14418 24670 14420 24722
rect 14140 24668 14420 24670
rect 14140 24388 14196 24668
rect 14364 24658 14420 24668
rect 14812 24612 14868 24622
rect 14812 24518 14868 24556
rect 13804 24332 14196 24388
rect 14252 24500 14308 24510
rect 12796 23998 12798 24050
rect 12850 23998 12852 24050
rect 12796 23986 12852 23998
rect 13692 24050 13748 24062
rect 13692 23998 13694 24050
rect 13746 23998 13748 24050
rect 13692 23940 13748 23998
rect 13692 23874 13748 23884
rect 12684 23774 12686 23826
rect 12738 23774 12740 23826
rect 12684 23762 12740 23774
rect 12908 23826 12964 23838
rect 12908 23774 12910 23826
rect 12962 23774 12964 23826
rect 12908 23380 12964 23774
rect 12908 23314 12964 23324
rect 13804 23268 13860 24332
rect 14140 24164 14196 24174
rect 13916 23380 13972 23390
rect 13916 23286 13972 23324
rect 13468 23266 13860 23268
rect 13468 23214 13806 23266
rect 13858 23214 13860 23266
rect 13468 23212 13860 23214
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 12908 21812 12964 21822
rect 9996 21700 10052 21710
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 4172 21410 4228 21420
rect 9996 21474 10052 21644
rect 12908 21586 12964 21756
rect 13468 21810 13524 23212
rect 13804 23202 13860 23212
rect 14140 23266 14196 24108
rect 14140 23214 14142 23266
rect 14194 23214 14196 23266
rect 14140 23202 14196 23214
rect 13468 21758 13470 21810
rect 13522 21758 13524 21810
rect 12908 21534 12910 21586
rect 12962 21534 12964 21586
rect 9996 21422 9998 21474
rect 10050 21422 10052 21474
rect 9996 21410 10052 21422
rect 12124 21474 12180 21486
rect 12124 21422 12126 21474
rect 12178 21422 12180 21474
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 9996 21140 10052 21150
rect 1932 20850 1988 20860
rect 2044 20914 2100 20926
rect 2044 20862 2046 20914
rect 2098 20862 2100 20914
rect 2044 20244 2100 20862
rect 9996 20914 10052 21084
rect 9996 20862 9998 20914
rect 10050 20862 10052 20914
rect 9996 20850 10052 20862
rect 12124 20916 12180 21422
rect 12124 20850 12180 20860
rect 4284 20804 4340 20814
rect 4284 20710 4340 20748
rect 12908 20802 12964 21534
rect 13244 21698 13300 21710
rect 13244 21646 13246 21698
rect 13298 21646 13300 21698
rect 13132 21364 13188 21374
rect 12908 20750 12910 20802
rect 12962 20750 12964 20802
rect 12908 20738 12964 20750
rect 13020 21362 13188 21364
rect 13020 21310 13134 21362
rect 13186 21310 13188 21362
rect 13020 21308 13188 21310
rect 12124 20692 12180 20702
rect 12124 20690 12404 20692
rect 12124 20638 12126 20690
rect 12178 20638 12404 20690
rect 12124 20636 12404 20638
rect 12124 20626 12180 20636
rect 2044 20178 2100 20188
rect 12348 20242 12404 20636
rect 12348 20190 12350 20242
rect 12402 20190 12404 20242
rect 12348 20178 12404 20190
rect 13020 20188 13076 21308
rect 13132 21298 13188 21308
rect 13244 21140 13300 21646
rect 13468 21364 13524 21758
rect 14140 21812 14196 21822
rect 14252 21812 14308 24444
rect 15148 24276 15204 25228
rect 15260 25282 15316 25294
rect 15260 25230 15262 25282
rect 15314 25230 15316 25282
rect 15260 25060 15316 25230
rect 16268 25284 16324 25294
rect 16268 25190 16324 25228
rect 16828 25284 16884 25454
rect 16828 25218 16884 25228
rect 15260 25004 16100 25060
rect 16044 24946 16100 25004
rect 16044 24894 16046 24946
rect 16098 24894 16100 24946
rect 16044 24882 16100 24894
rect 16156 24610 16212 24622
rect 16156 24558 16158 24610
rect 16210 24558 16212 24610
rect 15148 24220 15540 24276
rect 15484 23380 15540 24220
rect 16156 24164 16212 24558
rect 15932 24108 16156 24164
rect 15484 23266 15540 23324
rect 15820 23826 15876 23838
rect 15820 23774 15822 23826
rect 15874 23774 15876 23826
rect 15820 23378 15876 23774
rect 15820 23326 15822 23378
rect 15874 23326 15876 23378
rect 15820 23314 15876 23326
rect 15484 23214 15486 23266
rect 15538 23214 15540 23266
rect 15484 23202 15540 23214
rect 15708 23268 15764 23278
rect 15708 23174 15764 23212
rect 14364 23154 14420 23166
rect 14364 23102 14366 23154
rect 14418 23102 14420 23154
rect 14364 21924 14420 23102
rect 15932 22930 15988 24108
rect 16156 24070 16212 24108
rect 16940 24612 16996 26124
rect 17500 26180 17556 26190
rect 17500 26086 17556 26124
rect 17948 25396 18004 26238
rect 17948 25330 18004 25340
rect 18284 26290 18340 26302
rect 18284 26238 18286 26290
rect 18338 26238 18340 26290
rect 16940 24052 16996 24556
rect 17052 24052 17108 24062
rect 16604 24050 17108 24052
rect 16604 23998 17054 24050
rect 17106 23998 17108 24050
rect 16604 23996 17108 23998
rect 15932 22878 15934 22930
rect 15986 22878 15988 22930
rect 15932 22596 15988 22878
rect 14364 21858 14420 21868
rect 15484 22540 15988 22596
rect 16044 23940 16100 23950
rect 14196 21756 14308 21812
rect 15036 21812 15092 21822
rect 14140 21718 14196 21756
rect 13468 21298 13524 21308
rect 13580 21588 13636 21598
rect 13244 21074 13300 21084
rect 13356 20916 13412 20926
rect 13356 20580 13412 20860
rect 13468 20804 13524 20814
rect 13580 20804 13636 21532
rect 13468 20802 13636 20804
rect 13468 20750 13470 20802
rect 13522 20750 13636 20802
rect 13468 20748 13636 20750
rect 13692 21586 13748 21598
rect 13692 21534 13694 21586
rect 13746 21534 13748 21586
rect 13468 20738 13524 20748
rect 13580 20580 13636 20590
rect 13356 20578 13636 20580
rect 13356 20526 13582 20578
rect 13634 20526 13636 20578
rect 13356 20524 13636 20526
rect 13580 20514 13636 20524
rect 13692 20188 13748 21534
rect 14924 21588 14980 21598
rect 14924 21494 14980 21532
rect 14364 21364 14420 21374
rect 12572 20132 12628 20142
rect 12572 20038 12628 20076
rect 12684 20132 13076 20188
rect 13468 20132 13748 20188
rect 13804 20690 13860 20702
rect 13804 20638 13806 20690
rect 13858 20638 13860 20690
rect 12684 20130 12740 20132
rect 12684 20078 12686 20130
rect 12738 20078 12740 20130
rect 12684 20066 12740 20078
rect 4284 20020 4340 20030
rect 4284 19926 4340 19964
rect 13020 20020 13076 20030
rect 13020 19906 13076 19964
rect 13020 19854 13022 19906
rect 13074 19854 13076 19906
rect 13020 19842 13076 19854
rect 1932 19796 1988 19806
rect 1932 19702 1988 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 13468 18452 13524 20132
rect 12908 18396 13524 18452
rect 13804 19684 13860 20638
rect 14028 20692 14084 20702
rect 14028 20598 14084 20636
rect 14364 20690 14420 21308
rect 15036 20916 15092 21756
rect 15148 21700 15204 21710
rect 15148 21606 15204 21644
rect 15260 21586 15316 21598
rect 15260 21534 15262 21586
rect 15314 21534 15316 21586
rect 15260 21364 15316 21534
rect 15260 21298 15316 21308
rect 15148 20916 15204 20926
rect 15036 20860 15148 20916
rect 15148 20822 15204 20860
rect 14364 20638 14366 20690
rect 14418 20638 14420 20690
rect 14364 20626 14420 20638
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17778 1988 17790
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 16884 1988 17726
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 10332 17668 10388 17678
rect 1932 16818 1988 16828
rect 4284 16882 4340 16894
rect 4284 16830 4286 16882
rect 4338 16830 4340 16882
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4284 16324 4340 16830
rect 10332 16770 10388 17612
rect 12572 17668 12628 17678
rect 12572 17574 12628 17612
rect 12908 17666 12964 18396
rect 12908 17614 12910 17666
rect 12962 17614 12964 17666
rect 12908 17602 12964 17614
rect 12796 17556 12852 17566
rect 12796 17462 12852 17500
rect 12460 17444 12516 17454
rect 13244 17444 13300 18396
rect 13356 17668 13412 17678
rect 13356 17574 13412 17612
rect 13804 17666 13860 19628
rect 14700 20578 14756 20590
rect 14700 20526 14702 20578
rect 14754 20526 14756 20578
rect 14476 18452 14532 18462
rect 14700 18452 14756 20526
rect 15148 19906 15204 19918
rect 15148 19854 15150 19906
rect 15202 19854 15204 19906
rect 14924 19460 14980 19470
rect 15148 19460 15204 19854
rect 14924 19458 15204 19460
rect 14924 19406 14926 19458
rect 14978 19406 15204 19458
rect 14924 19404 15204 19406
rect 15260 19460 15316 19470
rect 15484 19460 15540 22540
rect 15932 22370 15988 22382
rect 15932 22318 15934 22370
rect 15986 22318 15988 22370
rect 15932 21924 15988 22318
rect 16044 22370 16100 23884
rect 16604 23938 16660 23996
rect 17052 23986 17108 23996
rect 16604 23886 16606 23938
rect 16658 23886 16660 23938
rect 16604 23874 16660 23886
rect 16828 23828 16884 23838
rect 16268 23154 16324 23166
rect 16268 23102 16270 23154
rect 16322 23102 16324 23154
rect 16268 22482 16324 23102
rect 16268 22430 16270 22482
rect 16322 22430 16324 22482
rect 16268 22418 16324 22430
rect 16044 22318 16046 22370
rect 16098 22318 16100 22370
rect 16044 22306 16100 22318
rect 16492 22370 16548 22382
rect 16492 22318 16494 22370
rect 16546 22318 16548 22370
rect 15932 21858 15988 21868
rect 15708 20916 15764 20926
rect 15764 20860 15876 20916
rect 15708 20822 15764 20860
rect 15820 20020 15876 20860
rect 16492 20132 16548 22318
rect 16268 20020 16324 20030
rect 15820 20018 16212 20020
rect 15820 19966 15822 20018
rect 15874 19966 16212 20018
rect 15820 19964 16212 19966
rect 15260 19458 15540 19460
rect 15260 19406 15262 19458
rect 15314 19406 15540 19458
rect 15260 19404 15540 19406
rect 15596 19796 15652 19806
rect 14924 19394 14980 19404
rect 15260 19394 15316 19404
rect 15036 19234 15092 19246
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 14700 18396 14868 18452
rect 14476 17780 14532 18396
rect 14028 17778 14532 17780
rect 14028 17726 14478 17778
rect 14530 17726 14532 17778
rect 14028 17724 14532 17726
rect 13804 17614 13806 17666
rect 13858 17614 13860 17666
rect 13804 17602 13860 17614
rect 13916 17666 13972 17678
rect 13916 17614 13918 17666
rect 13970 17614 13972 17666
rect 13580 17444 13636 17454
rect 13244 17388 13412 17444
rect 12460 16994 12516 17388
rect 12460 16942 12462 16994
rect 12514 16942 12516 16994
rect 12460 16930 12516 16942
rect 13244 16884 13300 16894
rect 13244 16790 13300 16828
rect 10332 16718 10334 16770
rect 10386 16718 10388 16770
rect 10332 16706 10388 16718
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4284 16258 4340 16268
rect 1932 16146 1988 16156
rect 9996 16210 10052 16222
rect 9996 16158 9998 16210
rect 10050 16158 10052 16210
rect 9996 16100 10052 16158
rect 13356 16212 13412 17388
rect 13580 17350 13636 17388
rect 9996 16034 10052 16044
rect 12908 16098 12964 16110
rect 12908 16046 12910 16098
rect 12962 16046 12964 16098
rect 12124 15988 12180 15998
rect 12124 15894 12180 15932
rect 12908 15540 12964 16046
rect 13356 16100 13412 16156
rect 13692 16884 13748 16894
rect 13468 16100 13524 16110
rect 13356 16098 13524 16100
rect 13356 16046 13470 16098
rect 13522 16046 13524 16098
rect 13356 16044 13524 16046
rect 13468 16034 13524 16044
rect 13132 15540 13188 15550
rect 13692 15540 13748 16828
rect 13916 16660 13972 17614
rect 14028 16884 14084 17724
rect 14476 17714 14532 17724
rect 14700 18228 14756 18238
rect 14700 16994 14756 18172
rect 14812 18116 14868 18396
rect 14812 18050 14868 18060
rect 15036 18340 15092 19182
rect 15484 19236 15540 19246
rect 15596 19236 15652 19740
rect 15484 19234 15652 19236
rect 15484 19182 15486 19234
rect 15538 19182 15652 19234
rect 15484 19180 15652 19182
rect 15484 19170 15540 19180
rect 15820 18452 15876 19964
rect 16156 19346 16212 19964
rect 16268 19926 16324 19964
rect 16268 19796 16324 19806
rect 16268 19702 16324 19740
rect 16492 19796 16548 20076
rect 16828 22146 16884 23772
rect 18284 23604 18340 26238
rect 18508 26292 18564 26302
rect 18956 26292 19012 26796
rect 18508 26198 18564 26236
rect 18620 26290 19012 26292
rect 18620 26238 18958 26290
rect 19010 26238 19012 26290
rect 18620 26236 19012 26238
rect 18620 26180 18676 26236
rect 18956 26226 19012 26236
rect 19292 26292 19348 26302
rect 19348 26236 19460 26292
rect 19292 26226 19348 26236
rect 18508 25620 18564 25630
rect 18620 25620 18676 26124
rect 18508 25618 18676 25620
rect 18508 25566 18510 25618
rect 18562 25566 18676 25618
rect 18508 25564 18676 25566
rect 19180 25732 19236 25742
rect 18508 25554 18564 25564
rect 17388 23380 17444 23390
rect 17388 23286 17444 23324
rect 18284 23268 18340 23548
rect 18284 23174 18340 23212
rect 18508 25396 18564 25406
rect 17612 23154 17668 23166
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 16828 22094 16830 22146
rect 16882 22094 16884 22146
rect 16604 19908 16660 19918
rect 16604 19814 16660 19852
rect 16492 19730 16548 19740
rect 16156 19294 16158 19346
rect 16210 19294 16212 19346
rect 16156 19282 16212 19294
rect 16828 19124 16884 22094
rect 17164 22370 17220 22382
rect 17164 22318 17166 22370
rect 17218 22318 17220 22370
rect 17164 21700 17220 22318
rect 17276 22372 17332 22382
rect 17276 22278 17332 22316
rect 17612 22372 17668 23102
rect 18172 22428 18452 22484
rect 17612 22306 17668 22316
rect 17948 22372 18004 22382
rect 18004 22316 18116 22372
rect 17948 22278 18004 22316
rect 18060 22036 18116 22316
rect 18172 22258 18228 22428
rect 18172 22206 18174 22258
rect 18226 22206 18228 22258
rect 18172 22194 18228 22206
rect 18284 22260 18340 22270
rect 18060 21980 18228 22036
rect 17948 21924 18004 21934
rect 17948 21810 18004 21868
rect 17948 21758 17950 21810
rect 18002 21758 18004 21810
rect 17948 21746 18004 21758
rect 17164 21644 17444 21700
rect 17388 21252 17444 21644
rect 17836 21586 17892 21598
rect 17836 21534 17838 21586
rect 17890 21534 17892 21586
rect 17500 21476 17556 21486
rect 17500 21382 17556 21420
rect 17836 21252 17892 21534
rect 18060 21476 18116 21486
rect 18060 21382 18116 21420
rect 17388 21196 17892 21252
rect 18060 21252 18116 21262
rect 16828 19058 16884 19068
rect 16380 19012 16436 19022
rect 15820 18386 15876 18396
rect 16044 18452 16100 18462
rect 16044 18450 16212 18452
rect 16044 18398 16046 18450
rect 16098 18398 16212 18450
rect 16044 18396 16212 18398
rect 16044 18386 16100 18396
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 14028 16790 14084 16828
rect 13916 16604 14084 16660
rect 13804 16100 13860 16110
rect 13804 16006 13860 16044
rect 14028 16100 14084 16604
rect 14028 16034 14084 16044
rect 14700 16100 14756 16110
rect 15036 16100 15092 18284
rect 16156 18340 16212 18396
rect 16380 18450 16436 18956
rect 16380 18398 16382 18450
rect 16434 18398 16436 18450
rect 16380 18386 16436 18398
rect 16940 19010 16996 19022
rect 16940 18958 16942 19010
rect 16994 18958 16996 19010
rect 16044 18228 16100 18238
rect 16044 18134 16100 18172
rect 16156 17892 16212 18284
rect 16156 17826 16212 17836
rect 16828 17556 16884 17566
rect 16828 16770 16884 17500
rect 16828 16718 16830 16770
rect 16882 16718 16884 16770
rect 16828 16706 16884 16718
rect 16940 16212 16996 18958
rect 17276 19010 17332 19022
rect 17276 18958 17278 19010
rect 17330 18958 17332 19010
rect 14700 16098 15092 16100
rect 14700 16046 14702 16098
rect 14754 16046 15092 16098
rect 14700 16044 15092 16046
rect 16380 16100 16436 16110
rect 14700 16034 14756 16044
rect 16380 16006 16436 16044
rect 16828 16100 16884 16110
rect 16940 16100 16996 16156
rect 16828 16098 16996 16100
rect 16828 16046 16830 16098
rect 16882 16046 16996 16098
rect 16828 16044 16996 16046
rect 17052 18452 17108 18462
rect 17052 17778 17108 18396
rect 17276 18452 17332 18958
rect 17612 18676 17668 21196
rect 18060 19234 18116 21196
rect 18172 19906 18228 21980
rect 18284 21586 18340 22204
rect 18284 21534 18286 21586
rect 18338 21534 18340 21586
rect 18284 21522 18340 21534
rect 18172 19854 18174 19906
rect 18226 19854 18228 19906
rect 18172 19842 18228 19854
rect 18396 19908 18452 22428
rect 18508 20692 18564 25340
rect 19068 25284 19124 25294
rect 18956 23938 19012 23950
rect 18956 23886 18958 23938
rect 19010 23886 19012 23938
rect 18956 23828 19012 23886
rect 18956 23762 19012 23772
rect 19068 23380 19124 25228
rect 19180 24162 19236 25676
rect 19404 25618 19460 26236
rect 19516 26180 19572 27134
rect 20412 27076 20468 27086
rect 21532 27076 21588 27086
rect 20412 27074 21252 27076
rect 20412 27022 20414 27074
rect 20466 27022 21252 27074
rect 20412 27020 21252 27022
rect 20412 27010 20468 27020
rect 19852 26964 19908 26974
rect 19852 26870 19908 26908
rect 20300 26964 20356 26974
rect 19740 26852 19796 26862
rect 19628 26850 19796 26852
rect 19628 26798 19742 26850
rect 19794 26798 19796 26850
rect 19628 26796 19796 26798
rect 19628 26402 19684 26796
rect 19740 26786 19796 26796
rect 20076 26852 20132 26862
rect 20076 26850 20244 26852
rect 20076 26798 20078 26850
rect 20130 26798 20244 26850
rect 20076 26796 20244 26798
rect 20076 26786 20132 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20188 26516 20244 26796
rect 19628 26350 19630 26402
rect 19682 26350 19684 26402
rect 19628 26338 19684 26350
rect 20076 26460 20244 26516
rect 19516 26124 19908 26180
rect 19404 25566 19406 25618
rect 19458 25566 19460 25618
rect 19404 25554 19460 25566
rect 19292 25506 19348 25518
rect 19292 25454 19294 25506
rect 19346 25454 19348 25506
rect 19292 25396 19348 25454
rect 19852 25506 19908 26124
rect 20076 25732 20132 26460
rect 20076 25666 20132 25676
rect 19852 25454 19854 25506
rect 19906 25454 19908 25506
rect 19852 25442 19908 25454
rect 19292 25330 19348 25340
rect 20188 25396 20244 25406
rect 19516 25282 19572 25294
rect 19740 25284 19796 25322
rect 19516 25230 19518 25282
rect 19570 25230 19572 25282
rect 19516 24724 19572 25230
rect 19516 24658 19572 24668
rect 19628 25228 19740 25284
rect 19628 24500 19684 25228
rect 19740 25218 19796 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19852 24948 19908 24958
rect 19852 24854 19908 24892
rect 20188 24946 20244 25340
rect 20188 24894 20190 24946
rect 20242 24894 20244 24946
rect 20188 24882 20244 24894
rect 20300 24948 20356 26908
rect 20748 26852 20804 26862
rect 20748 26758 20804 26796
rect 21196 25506 21252 27020
rect 21532 26982 21588 27020
rect 21756 26178 21812 37998
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24556 31948 24612 37998
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 40236 36372 40292 36382
rect 40236 36278 40292 36316
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 24332 31892 24612 31948
rect 24332 27186 24388 31892
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 24332 27134 24334 27186
rect 24386 27134 24388 27186
rect 24108 27076 24164 27086
rect 22204 26964 22260 26974
rect 21980 26962 22260 26964
rect 21980 26910 22206 26962
rect 22258 26910 22260 26962
rect 21980 26908 22260 26910
rect 24108 26908 24164 27020
rect 21980 26514 22036 26908
rect 22204 26898 22260 26908
rect 23996 26852 24164 26908
rect 21980 26462 21982 26514
rect 22034 26462 22036 26514
rect 21980 26450 22036 26462
rect 22204 26740 22260 26750
rect 22204 26514 22260 26684
rect 22988 26516 23044 26526
rect 22204 26462 22206 26514
rect 22258 26462 22260 26514
rect 22204 26450 22260 26462
rect 22316 26514 23044 26516
rect 22316 26462 22990 26514
rect 23042 26462 23044 26514
rect 22316 26460 23044 26462
rect 22316 26402 22372 26460
rect 22988 26450 23044 26460
rect 22316 26350 22318 26402
rect 22370 26350 22372 26402
rect 22316 26338 22372 26350
rect 21756 26126 21758 26178
rect 21810 26126 21812 26178
rect 21756 26068 21812 26126
rect 21196 25454 21198 25506
rect 21250 25454 21252 25506
rect 21196 25442 21252 25454
rect 21420 26012 21812 26068
rect 22652 26290 22708 26302
rect 22652 26238 22654 26290
rect 22706 26238 22708 26290
rect 21420 25394 21476 26012
rect 21420 25342 21422 25394
rect 21474 25342 21476 25394
rect 21420 25330 21476 25342
rect 21532 25394 21588 25406
rect 21532 25342 21534 25394
rect 21586 25342 21588 25394
rect 21532 25284 21588 25342
rect 21532 25218 21588 25228
rect 22652 25284 22708 26238
rect 22876 26292 22932 26302
rect 22876 26198 22932 26236
rect 23100 26290 23156 26302
rect 23100 26238 23102 26290
rect 23154 26238 23156 26290
rect 22652 25218 22708 25228
rect 20300 24882 20356 24892
rect 21308 24834 21364 24846
rect 21308 24782 21310 24834
rect 21362 24782 21364 24834
rect 19404 24444 19684 24500
rect 19740 24722 19796 24734
rect 19740 24670 19742 24722
rect 19794 24670 19796 24722
rect 19180 24110 19182 24162
rect 19234 24110 19236 24162
rect 19180 24098 19236 24110
rect 19292 24276 19348 24286
rect 18620 23154 18676 23166
rect 18620 23102 18622 23154
rect 18674 23102 18676 23154
rect 18620 22260 18676 23102
rect 19068 22482 19124 23324
rect 19180 23716 19236 23726
rect 19180 23154 19236 23660
rect 19292 23714 19348 24220
rect 19292 23662 19294 23714
rect 19346 23662 19348 23714
rect 19292 23604 19348 23662
rect 19292 23538 19348 23548
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 19180 23090 19236 23102
rect 19068 22430 19070 22482
rect 19122 22430 19124 22482
rect 19068 22418 19124 22430
rect 19404 22482 19460 24444
rect 19740 24276 19796 24670
rect 19964 24724 20020 24734
rect 19964 24630 20020 24668
rect 21308 24724 21364 24782
rect 19740 24210 19796 24220
rect 19516 23828 19572 23838
rect 19516 23714 19572 23772
rect 20748 23826 20804 23838
rect 20748 23774 20750 23826
rect 20802 23774 20804 23826
rect 19516 23662 19518 23714
rect 19570 23662 19572 23714
rect 19516 22596 19572 23662
rect 20412 23714 20468 23726
rect 20412 23662 20414 23714
rect 20466 23662 20468 23714
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19964 23042 20020 23054
rect 19964 22990 19966 23042
rect 20018 22990 20020 23042
rect 19516 22540 19684 22596
rect 19404 22430 19406 22482
rect 19458 22430 19460 22482
rect 19404 22418 19460 22430
rect 19292 22372 19348 22382
rect 18732 22260 18788 22270
rect 18620 22258 18788 22260
rect 18620 22206 18734 22258
rect 18786 22206 18788 22258
rect 18620 22204 18788 22206
rect 18732 21588 18788 22204
rect 19292 22258 19348 22316
rect 19292 22206 19294 22258
rect 19346 22206 19348 22258
rect 19292 22194 19348 22206
rect 19516 22370 19572 22382
rect 19516 22318 19518 22370
rect 19570 22318 19572 22370
rect 19068 21812 19124 21822
rect 19068 21718 19124 21756
rect 18844 21588 18900 21598
rect 18732 21586 18900 21588
rect 18732 21534 18846 21586
rect 18898 21534 18900 21586
rect 18732 21532 18900 21534
rect 18844 21476 18900 21532
rect 19404 21588 19460 21598
rect 19404 21494 19460 21532
rect 18844 21410 18900 21420
rect 18620 20692 18676 20702
rect 18508 20636 18620 20692
rect 18620 20626 18676 20636
rect 19404 20692 19460 20702
rect 18956 20242 19012 20254
rect 18956 20190 18958 20242
rect 19010 20190 19012 20242
rect 18956 20188 19012 20190
rect 18060 19182 18062 19234
rect 18114 19182 18116 19234
rect 18060 19170 18116 19182
rect 17724 19124 17780 19134
rect 17724 19030 17780 19068
rect 17836 19012 17892 19022
rect 17836 18918 17892 18956
rect 17724 18676 17780 18686
rect 17612 18674 18004 18676
rect 17612 18622 17726 18674
rect 17778 18622 18004 18674
rect 17612 18620 18004 18622
rect 17724 18610 17780 18620
rect 17276 18386 17332 18396
rect 17500 18452 17556 18462
rect 17500 18450 17668 18452
rect 17500 18398 17502 18450
rect 17554 18398 17668 18450
rect 17500 18396 17668 18398
rect 17500 18386 17556 18396
rect 17052 17726 17054 17778
rect 17106 17726 17108 17778
rect 16828 16034 16884 16044
rect 14364 15988 14420 15998
rect 14140 15986 14420 15988
rect 14140 15934 14366 15986
rect 14418 15934 14420 15986
rect 14140 15932 14420 15934
rect 13916 15874 13972 15886
rect 13916 15822 13918 15874
rect 13970 15822 13972 15874
rect 13916 15652 13972 15822
rect 14140 15652 14196 15932
rect 14364 15922 14420 15932
rect 14476 15988 14532 15998
rect 14476 15894 14532 15932
rect 13916 15596 14196 15652
rect 16492 15874 16548 15886
rect 16492 15822 16494 15874
rect 16546 15822 16548 15874
rect 12908 15538 13748 15540
rect 12908 15486 13134 15538
rect 13186 15486 13748 15538
rect 12908 15484 13748 15486
rect 13132 15474 13188 15484
rect 13692 15316 13748 15484
rect 13916 15316 13972 15326
rect 13692 15314 13972 15316
rect 13692 15262 13918 15314
rect 13970 15262 13972 15314
rect 13692 15260 13972 15262
rect 13916 15250 13972 15260
rect 14700 15202 14756 15214
rect 14700 15150 14702 15202
rect 14754 15150 14756 15202
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14700 14756 14756 15150
rect 16492 15092 16548 15822
rect 16604 15874 16660 15886
rect 16604 15822 16606 15874
rect 16658 15822 16660 15874
rect 16604 15148 16660 15822
rect 17052 15876 17108 17726
rect 17612 18116 17668 18396
rect 17612 17668 17668 18060
rect 17724 17668 17780 17678
rect 17612 17612 17724 17668
rect 17948 17668 18004 18620
rect 18284 18340 18340 18350
rect 18396 18340 18452 19852
rect 18508 20132 19012 20188
rect 18508 20020 18564 20132
rect 18508 19796 18564 19964
rect 18620 20020 18676 20030
rect 18620 20018 19012 20020
rect 18620 19966 18622 20018
rect 18674 19966 19012 20018
rect 18620 19964 19012 19966
rect 18620 19954 18676 19964
rect 18956 19908 19012 19964
rect 19180 20018 19236 20030
rect 19180 19966 19182 20018
rect 19234 19966 19236 20018
rect 19180 19908 19236 19966
rect 18956 19852 19236 19908
rect 18844 19796 18900 19806
rect 18508 19740 18788 19796
rect 18508 19236 18564 19246
rect 18508 19234 18676 19236
rect 18508 19182 18510 19234
rect 18562 19182 18676 19234
rect 18508 19180 18676 19182
rect 18508 19170 18564 19180
rect 18620 18676 18676 19180
rect 18732 19122 18788 19740
rect 18844 19702 18900 19740
rect 18732 19070 18734 19122
rect 18786 19070 18788 19122
rect 18732 19058 18788 19070
rect 19180 19234 19236 19852
rect 19404 19572 19460 20636
rect 19516 20132 19572 22318
rect 19628 22148 19684 22540
rect 19964 22148 20020 22990
rect 19628 22092 20020 22148
rect 20300 22370 20356 22382
rect 20300 22318 20302 22370
rect 20354 22318 20356 22370
rect 19628 20132 19684 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 21822
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19964 20244 20020 20254
rect 20188 20244 20244 21756
rect 19964 20242 20244 20244
rect 19964 20190 19966 20242
rect 20018 20190 20244 20242
rect 19964 20188 20244 20190
rect 19964 20178 20020 20188
rect 19740 20132 19796 20142
rect 19628 20130 19908 20132
rect 19628 20078 19742 20130
rect 19794 20078 19908 20130
rect 19628 20076 19908 20078
rect 19516 20018 19572 20076
rect 19740 20066 19796 20076
rect 19516 19966 19518 20018
rect 19570 19966 19572 20018
rect 19516 19954 19572 19966
rect 19628 19796 19684 19806
rect 19628 19702 19684 19740
rect 19404 19516 19796 19572
rect 19180 19182 19182 19234
rect 19234 19182 19236 19234
rect 19180 18788 19236 19182
rect 19516 19236 19572 19246
rect 19404 19012 19460 19022
rect 19516 19012 19572 19180
rect 19740 19122 19796 19516
rect 19740 19070 19742 19122
rect 19794 19070 19796 19122
rect 19740 19058 19796 19070
rect 19404 19010 19572 19012
rect 19404 18958 19406 19010
rect 19458 18958 19572 19010
rect 19404 18956 19572 18958
rect 19852 19012 19908 20076
rect 20188 20018 20244 20030
rect 20188 19966 20190 20018
rect 20242 19966 20244 20018
rect 20188 19236 20244 19966
rect 20300 20020 20356 22318
rect 20412 22148 20468 23662
rect 20636 23714 20692 23726
rect 20636 23662 20638 23714
rect 20690 23662 20692 23714
rect 20636 23604 20692 23662
rect 20636 23538 20692 23548
rect 20412 22082 20468 22092
rect 20748 21812 20804 23774
rect 21308 23604 21364 24668
rect 21644 24722 21700 24734
rect 21644 24670 21646 24722
rect 21698 24670 21700 24722
rect 21532 23604 21588 23614
rect 21308 23548 21532 23604
rect 21308 22260 21364 22270
rect 21308 22166 21364 22204
rect 20748 21746 20804 21756
rect 21196 21812 21252 21822
rect 20300 19954 20356 19964
rect 20412 21476 20468 21486
rect 20188 19170 20244 19180
rect 20412 19122 20468 21420
rect 20412 19070 20414 19122
rect 20466 19070 20468 19122
rect 20412 19058 20468 19070
rect 20524 20356 20580 20366
rect 19964 19012 20020 19022
rect 19852 18956 19964 19012
rect 19404 18946 19460 18956
rect 19180 18732 19460 18788
rect 18620 18620 19348 18676
rect 18620 18450 18676 18620
rect 18620 18398 18622 18450
rect 18674 18398 18676 18450
rect 18620 18386 18676 18398
rect 18284 18338 18452 18340
rect 18284 18286 18286 18338
rect 18338 18286 18452 18338
rect 18284 18284 18452 18286
rect 18284 18004 18340 18284
rect 18284 17938 18340 17948
rect 18060 17892 18116 17902
rect 18060 17798 18116 17836
rect 18844 17890 18900 18620
rect 19068 18452 19124 18462
rect 19068 18116 19124 18396
rect 19292 18450 19348 18620
rect 19292 18398 19294 18450
rect 19346 18398 19348 18450
rect 19292 18386 19348 18398
rect 19068 18050 19124 18060
rect 18844 17838 18846 17890
rect 18898 17838 18900 17890
rect 18060 17668 18116 17678
rect 17948 17666 18228 17668
rect 17948 17614 18062 17666
rect 18114 17614 18228 17666
rect 17948 17612 18228 17614
rect 17388 17556 17444 17566
rect 17388 17462 17444 17500
rect 17724 17554 17780 17612
rect 18060 17602 18116 17612
rect 17724 17502 17726 17554
rect 17778 17502 17780 17554
rect 17724 17490 17780 17502
rect 18172 16994 18228 17612
rect 18172 16942 18174 16994
rect 18226 16942 18228 16994
rect 18172 16930 18228 16942
rect 18396 17554 18452 17566
rect 18396 17502 18398 17554
rect 18450 17502 18452 17554
rect 18396 16996 18452 17502
rect 18732 17556 18788 17566
rect 18732 17462 18788 17500
rect 18844 17106 18900 17838
rect 19404 17892 19460 18732
rect 19404 17826 19460 17836
rect 18844 17054 18846 17106
rect 18898 17054 18900 17106
rect 18844 17042 18900 17054
rect 19516 17108 19572 18956
rect 19964 18946 20020 18956
rect 20076 19012 20132 19022
rect 20076 19010 20244 19012
rect 20076 18958 20078 19010
rect 20130 18958 20244 19010
rect 20076 18956 20244 18958
rect 20076 18946 20132 18956
rect 20188 18900 20244 18956
rect 20524 18900 20580 20300
rect 20860 20132 20916 20142
rect 20748 19236 20804 19246
rect 20748 19142 20804 19180
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18844 20580 18900
rect 20188 18676 20244 18844
rect 19852 18620 20244 18676
rect 20748 18676 20804 18686
rect 20860 18676 20916 20076
rect 20748 18674 20916 18676
rect 20748 18622 20750 18674
rect 20802 18622 20916 18674
rect 20748 18620 20916 18622
rect 20972 19236 21028 19246
rect 19852 18340 19908 18620
rect 20748 18610 20804 18620
rect 19852 18246 19908 18284
rect 20188 18338 20244 18350
rect 20188 18286 20190 18338
rect 20242 18286 20244 18338
rect 20188 18228 20244 18286
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 20188 17108 20244 18172
rect 20636 17892 20692 17902
rect 20636 17798 20692 17836
rect 20748 17556 20804 17566
rect 20748 17462 20804 17500
rect 19516 17052 19852 17108
rect 18396 16930 18452 16940
rect 18508 16994 18564 17006
rect 18508 16942 18510 16994
rect 18562 16942 18564 16994
rect 17948 16884 18004 16894
rect 17948 16790 18004 16828
rect 18508 16772 18564 16942
rect 19404 16996 19460 17006
rect 19180 16884 19236 16922
rect 19180 16818 19236 16828
rect 19404 16772 19460 16940
rect 19852 16994 19908 17052
rect 20076 17052 20244 17108
rect 19852 16942 19854 16994
rect 19906 16942 19908 16994
rect 19852 16930 19908 16942
rect 19964 16994 20020 17006
rect 19964 16942 19966 16994
rect 20018 16942 20020 16994
rect 19516 16772 19572 16782
rect 19404 16770 19572 16772
rect 19404 16718 19518 16770
rect 19570 16718 19572 16770
rect 19404 16716 19572 16718
rect 17612 16658 17668 16670
rect 17612 16606 17614 16658
rect 17666 16606 17668 16658
rect 17612 16324 17668 16606
rect 17164 16268 17668 16324
rect 17164 16098 17220 16268
rect 17164 16046 17166 16098
rect 17218 16046 17220 16098
rect 17164 16034 17220 16046
rect 18508 16100 18564 16716
rect 19516 16706 19572 16716
rect 19964 16772 20020 16942
rect 20076 16884 20132 17052
rect 20076 16818 20132 16828
rect 20188 16884 20244 16894
rect 20636 16884 20692 16894
rect 20188 16882 20692 16884
rect 20188 16830 20190 16882
rect 20242 16830 20638 16882
rect 20690 16830 20692 16882
rect 20188 16828 20692 16830
rect 20188 16818 20244 16828
rect 20636 16818 20692 16828
rect 19964 16706 20020 16716
rect 20860 16770 20916 16782
rect 20860 16718 20862 16770
rect 20914 16718 20916 16770
rect 18508 16034 18564 16044
rect 19180 16658 19236 16670
rect 19180 16606 19182 16658
rect 19234 16606 19236 16658
rect 17052 15820 17556 15876
rect 17500 15538 17556 15820
rect 17500 15486 17502 15538
rect 17554 15486 17556 15538
rect 16828 15202 16884 15214
rect 16828 15150 16830 15202
rect 16882 15150 16884 15202
rect 16828 15148 16884 15150
rect 16604 15092 16884 15148
rect 15820 15036 16548 15092
rect 14700 14690 14756 14700
rect 15708 14756 15764 14766
rect 15708 14662 15764 14700
rect 15820 14642 15876 15036
rect 15820 14590 15822 14642
rect 15874 14590 15876 14642
rect 15820 14578 15876 14590
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16828 8428 16884 15092
rect 17500 14532 17556 15486
rect 19180 15148 19236 16606
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20748 15428 20804 15438
rect 20860 15428 20916 16718
rect 20748 15426 20916 15428
rect 20748 15374 20750 15426
rect 20802 15374 20916 15426
rect 20748 15372 20916 15374
rect 20748 15362 20804 15372
rect 20076 15316 20132 15326
rect 20076 15222 20132 15260
rect 18620 15092 19236 15148
rect 18620 14642 18676 15092
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 20748 14644 20804 14654
rect 20972 14644 21028 19180
rect 21196 18562 21252 21756
rect 21308 20802 21364 20814
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 21308 20356 21364 20750
rect 21532 20690 21588 23548
rect 21644 23044 21700 24670
rect 21868 24052 21924 24062
rect 21868 24050 22260 24052
rect 21868 23998 21870 24050
rect 21922 23998 22260 24050
rect 21868 23996 22260 23998
rect 21868 23986 21924 23996
rect 22204 23940 22260 23996
rect 22652 23940 22708 23950
rect 22204 23938 22708 23940
rect 22204 23886 22654 23938
rect 22706 23886 22708 23938
rect 22204 23884 22708 23886
rect 22092 23826 22148 23838
rect 22092 23774 22094 23826
rect 22146 23774 22148 23826
rect 22092 23044 22148 23774
rect 21644 23042 22148 23044
rect 21644 22990 22094 23042
rect 22146 22990 22148 23042
rect 21644 22988 22148 22990
rect 21532 20638 21534 20690
rect 21586 20638 21588 20690
rect 21532 20626 21588 20638
rect 21308 20290 21364 20300
rect 21308 20132 21364 20142
rect 21308 19906 21364 20076
rect 21420 20020 21476 20030
rect 21756 20020 21812 22988
rect 22092 22978 22148 22988
rect 22204 23156 22260 23884
rect 22652 23874 22708 23884
rect 22764 23828 22820 23838
rect 22428 23716 22484 23726
rect 22764 23716 22820 23772
rect 22428 23714 22820 23716
rect 22428 23662 22430 23714
rect 22482 23662 22820 23714
rect 22428 23660 22820 23662
rect 22428 23650 22484 23660
rect 23100 23492 23156 26238
rect 23324 26290 23380 26302
rect 23324 26238 23326 26290
rect 23378 26238 23380 26290
rect 23324 25284 23380 26238
rect 23324 25218 23380 25228
rect 23996 25506 24052 26852
rect 24332 26292 24388 27134
rect 24780 27076 24836 27086
rect 24780 26982 24836 27020
rect 40236 26850 40292 26862
rect 40236 26798 40238 26850
rect 40290 26798 40292 26850
rect 24332 26226 24388 26236
rect 37884 26290 37940 26302
rect 37884 26238 37886 26290
rect 37938 26238 37940 26290
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 23996 25454 23998 25506
rect 24050 25454 24052 25506
rect 23212 23716 23268 23726
rect 23212 23622 23268 23660
rect 23996 23716 24052 25454
rect 26908 25620 26964 25630
rect 24780 25396 24836 25406
rect 24332 25394 24836 25396
rect 24332 25342 24782 25394
rect 24834 25342 24836 25394
rect 24332 25340 24836 25342
rect 24108 24164 24164 24174
rect 24108 23938 24164 24108
rect 24332 24050 24388 25340
rect 24780 25330 24836 25340
rect 25340 25284 25396 25294
rect 24332 23998 24334 24050
rect 24386 23998 24388 24050
rect 24332 23986 24388 23998
rect 24668 24500 24724 24510
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 24108 23874 24164 23886
rect 24668 23938 24724 24444
rect 25004 24164 25060 24174
rect 25060 24108 25172 24164
rect 25004 24098 25060 24108
rect 24668 23886 24670 23938
rect 24722 23886 24724 23938
rect 24668 23874 24724 23886
rect 25004 23938 25060 23950
rect 25004 23886 25006 23938
rect 25058 23886 25060 23938
rect 24220 23716 24276 23726
rect 24444 23716 24500 23726
rect 23996 23650 24052 23660
rect 24108 23714 24276 23716
rect 24108 23662 24222 23714
rect 24274 23662 24276 23714
rect 24108 23660 24276 23662
rect 23100 23426 23156 23436
rect 23884 23268 23940 23278
rect 24108 23268 24164 23660
rect 24220 23650 24276 23660
rect 24332 23714 24500 23716
rect 24332 23662 24446 23714
rect 24498 23662 24500 23714
rect 24332 23660 24500 23662
rect 23884 23266 24276 23268
rect 23884 23214 23886 23266
rect 23938 23214 24276 23266
rect 23884 23212 24276 23214
rect 23884 23202 23940 23212
rect 22092 22260 22148 22270
rect 22204 22260 22260 23100
rect 23100 23154 23156 23166
rect 23100 23102 23102 23154
rect 23154 23102 23156 23154
rect 22148 22204 22260 22260
rect 22428 23042 22484 23054
rect 22428 22990 22430 23042
rect 22482 22990 22484 23042
rect 22092 22194 22148 22204
rect 22316 21812 22372 21822
rect 21980 20916 22036 20926
rect 21980 20822 22036 20860
rect 22316 20802 22372 21756
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 22316 20738 22372 20750
rect 22428 20132 22484 22990
rect 22764 23044 22820 23054
rect 23100 23044 23156 23102
rect 23324 23156 23380 23166
rect 23324 23062 23380 23100
rect 22764 23042 23156 23044
rect 22764 22990 22766 23042
rect 22818 22990 23156 23042
rect 22764 22988 23156 22990
rect 22764 22978 22820 22988
rect 23100 22370 23156 22988
rect 23100 22318 23102 22370
rect 23154 22318 23156 22370
rect 22876 21924 22932 21934
rect 22876 20802 22932 21868
rect 23100 21700 23156 22318
rect 23548 22372 23604 22382
rect 23548 22370 24052 22372
rect 23548 22318 23550 22370
rect 23602 22318 24052 22370
rect 23548 22316 24052 22318
rect 23548 22306 23604 22316
rect 23100 21634 23156 21644
rect 22876 20750 22878 20802
rect 22930 20750 22932 20802
rect 22876 20244 22932 20750
rect 23324 21474 23380 21486
rect 23324 21422 23326 21474
rect 23378 21422 23380 21474
rect 23324 20804 23380 21422
rect 23324 20710 23380 20748
rect 23100 20244 23156 20254
rect 22876 20242 23156 20244
rect 22876 20190 23102 20242
rect 23154 20190 23156 20242
rect 22876 20188 23156 20190
rect 23100 20178 23156 20188
rect 22428 20066 22484 20076
rect 21420 20018 21812 20020
rect 21420 19966 21422 20018
rect 21474 19966 21812 20018
rect 21420 19964 21812 19966
rect 21868 20020 21924 20030
rect 21420 19954 21476 19964
rect 21308 19854 21310 19906
rect 21362 19854 21364 19906
rect 21308 19236 21364 19854
rect 21532 19236 21588 19246
rect 21364 19234 21588 19236
rect 21364 19182 21534 19234
rect 21586 19182 21588 19234
rect 21364 19180 21588 19182
rect 21308 19142 21364 19180
rect 21532 19170 21588 19180
rect 21644 19122 21700 19964
rect 21868 19348 21924 19964
rect 22540 20020 22596 20030
rect 22540 19926 22596 19964
rect 22764 20018 22820 20030
rect 22764 19966 22766 20018
rect 22818 19966 22820 20018
rect 22764 19908 22820 19966
rect 23772 20020 23828 20030
rect 23772 19926 23828 19964
rect 22764 19842 22820 19852
rect 23548 19908 23604 19918
rect 23548 19814 23604 19852
rect 21644 19070 21646 19122
rect 21698 19070 21700 19122
rect 21644 19058 21700 19070
rect 21756 19346 21924 19348
rect 21756 19294 21870 19346
rect 21922 19294 21924 19346
rect 21756 19292 21924 19294
rect 21308 19012 21364 19022
rect 21308 18674 21364 18956
rect 21308 18622 21310 18674
rect 21362 18622 21364 18674
rect 21308 18610 21364 18622
rect 21196 18510 21198 18562
rect 21250 18510 21252 18562
rect 21196 18498 21252 18510
rect 21532 18452 21588 18462
rect 21532 18358 21588 18396
rect 21084 16996 21140 17006
rect 21084 16902 21140 16940
rect 21308 16996 21364 17006
rect 21756 16996 21812 19292
rect 21868 19282 21924 19292
rect 22540 19234 22596 19246
rect 22540 19182 22542 19234
rect 22594 19182 22596 19234
rect 21980 19124 22036 19134
rect 21980 18562 22036 19068
rect 21980 18510 21982 18562
rect 22034 18510 22036 18562
rect 21980 18498 22036 18510
rect 22316 18452 22372 18462
rect 22316 18358 22372 18396
rect 22204 18116 22260 18126
rect 22204 17554 22260 18060
rect 22204 17502 22206 17554
rect 22258 17502 22260 17554
rect 22204 17490 22260 17502
rect 22540 17556 22596 19182
rect 23772 19234 23828 19246
rect 23772 19182 23774 19234
rect 23826 19182 23828 19234
rect 23212 18564 23268 18574
rect 22764 18450 22820 18462
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 22764 18228 22820 18398
rect 22764 18162 22820 18172
rect 22988 18452 23044 18462
rect 22988 17668 23044 18396
rect 22988 17574 23044 17612
rect 21308 16994 21812 16996
rect 21308 16942 21310 16994
rect 21362 16942 21812 16994
rect 21308 16940 21812 16942
rect 22540 17442 22596 17500
rect 23212 17554 23268 18508
rect 23324 18450 23380 18462
rect 23324 18398 23326 18450
rect 23378 18398 23380 18450
rect 23324 18340 23380 18398
rect 23772 18452 23828 19182
rect 23884 18564 23940 18574
rect 23884 18470 23940 18508
rect 23772 18386 23828 18396
rect 23660 18340 23716 18350
rect 23324 18274 23380 18284
rect 23436 18338 23716 18340
rect 23436 18286 23662 18338
rect 23714 18286 23716 18338
rect 23436 18284 23716 18286
rect 23212 17502 23214 17554
rect 23266 17502 23268 17554
rect 23212 17490 23268 17502
rect 22540 17390 22542 17442
rect 22594 17390 22596 17442
rect 21308 16930 21364 16940
rect 22540 15204 22596 17390
rect 23436 16770 23492 18284
rect 23660 18274 23716 18284
rect 23772 18228 23828 18238
rect 23772 17778 23828 18172
rect 23772 17726 23774 17778
rect 23826 17726 23828 17778
rect 23772 17714 23828 17726
rect 23996 18004 24052 22316
rect 24108 19796 24164 19806
rect 24108 19702 24164 19740
rect 24108 19234 24164 19246
rect 24108 19182 24110 19234
rect 24162 19182 24164 19234
rect 24108 18116 24164 19182
rect 24108 18050 24164 18060
rect 23996 17668 24052 17948
rect 24108 17668 24164 17678
rect 23996 17666 24164 17668
rect 23996 17614 24110 17666
rect 24162 17614 24164 17666
rect 23996 17612 24164 17614
rect 24108 17602 24164 17612
rect 23772 17108 23828 17118
rect 23772 16882 23828 17052
rect 24220 16996 24276 23212
rect 24332 21924 24388 23660
rect 24444 23650 24500 23660
rect 25004 23716 25060 23886
rect 25004 23650 25060 23660
rect 24556 22260 24612 22270
rect 24556 22258 24948 22260
rect 24556 22206 24558 22258
rect 24610 22206 24948 22258
rect 24556 22204 24948 22206
rect 24556 22194 24612 22204
rect 24444 22148 24500 22158
rect 24444 22036 24500 22092
rect 24444 21980 24612 22036
rect 24332 21858 24388 21868
rect 24444 21812 24500 21822
rect 24444 20130 24500 21756
rect 24444 20078 24446 20130
rect 24498 20078 24500 20130
rect 24332 19348 24388 19358
rect 24444 19348 24500 20078
rect 24556 20130 24612 21980
rect 24556 20078 24558 20130
rect 24610 20078 24612 20130
rect 24556 20066 24612 20078
rect 24780 21588 24836 21598
rect 24780 20130 24836 21532
rect 24780 20078 24782 20130
rect 24834 20078 24836 20130
rect 24780 20066 24836 20078
rect 24892 20020 24948 22204
rect 25004 22148 25060 22158
rect 25004 22054 25060 22092
rect 25116 21812 25172 24108
rect 25228 23154 25284 23166
rect 25228 23102 25230 23154
rect 25282 23102 25284 23154
rect 25228 22148 25284 23102
rect 25228 22082 25284 22092
rect 25228 21812 25284 21822
rect 25116 21810 25284 21812
rect 25116 21758 25230 21810
rect 25282 21758 25284 21810
rect 25116 21756 25284 21758
rect 25228 21746 25284 21756
rect 25340 20130 25396 25228
rect 25564 24836 25620 24846
rect 25564 24742 25620 24780
rect 26908 24836 26964 25564
rect 27356 25620 27412 25630
rect 27356 25506 27412 25564
rect 27356 25454 27358 25506
rect 27410 25454 27412 25506
rect 27356 25442 27412 25454
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 27580 25284 27636 25294
rect 27580 25190 27636 25228
rect 28028 25282 28084 25294
rect 28028 25230 28030 25282
rect 28082 25230 28084 25282
rect 26908 24770 26964 24780
rect 25452 24500 25508 24510
rect 25452 24406 25508 24444
rect 26908 24052 26964 24062
rect 25788 23828 25844 23838
rect 25676 23826 25844 23828
rect 25676 23774 25790 23826
rect 25842 23774 25844 23826
rect 25676 23772 25844 23774
rect 25452 23492 25508 23502
rect 25452 23266 25508 23436
rect 25676 23378 25732 23772
rect 25788 23762 25844 23772
rect 25676 23326 25678 23378
rect 25730 23326 25732 23378
rect 25676 23314 25732 23326
rect 25452 23214 25454 23266
rect 25506 23214 25508 23266
rect 25452 23202 25508 23214
rect 25788 23154 25844 23166
rect 25788 23102 25790 23154
rect 25842 23102 25844 23154
rect 25788 22482 25844 23102
rect 25788 22430 25790 22482
rect 25842 22430 25844 22482
rect 25788 22418 25844 22430
rect 26124 23156 26180 23166
rect 26124 22370 26180 23100
rect 26124 22318 26126 22370
rect 26178 22318 26180 22370
rect 26124 22306 26180 22318
rect 25676 22260 25732 22270
rect 25676 22166 25732 22204
rect 25564 22146 25620 22158
rect 25564 22094 25566 22146
rect 25618 22094 25620 22146
rect 25564 21812 25620 22094
rect 25900 22146 25956 22158
rect 25900 22094 25902 22146
rect 25954 22094 25956 22146
rect 25900 21924 25956 22094
rect 25900 21858 25956 21868
rect 25564 21718 25620 21756
rect 25340 20078 25342 20130
rect 25394 20078 25396 20130
rect 25340 20066 25396 20078
rect 25452 21700 25508 21710
rect 25116 20020 25172 20030
rect 24892 20018 25172 20020
rect 24892 19966 25118 20018
rect 25170 19966 25172 20018
rect 24892 19964 25172 19966
rect 24332 19346 24500 19348
rect 24332 19294 24334 19346
rect 24386 19294 24500 19346
rect 24332 19292 24500 19294
rect 25116 19346 25172 19964
rect 25452 20018 25508 21644
rect 26012 21586 26068 21598
rect 26012 21534 26014 21586
rect 26066 21534 26068 21586
rect 26012 20916 26068 21534
rect 26236 21588 26292 21598
rect 26236 21494 26292 21532
rect 26572 21586 26628 21598
rect 26572 21534 26574 21586
rect 26626 21534 26628 21586
rect 26012 20850 26068 20860
rect 26460 21474 26516 21486
rect 26460 21422 26462 21474
rect 26514 21422 26516 21474
rect 26460 20132 26516 21422
rect 26460 20066 26516 20076
rect 25452 19966 25454 20018
rect 25506 19966 25508 20018
rect 25452 19954 25508 19966
rect 25788 20020 25844 20030
rect 25788 20018 25956 20020
rect 25788 19966 25790 20018
rect 25842 19966 25956 20018
rect 25788 19964 25956 19966
rect 25788 19954 25844 19964
rect 25116 19294 25118 19346
rect 25170 19294 25172 19346
rect 24332 19282 24388 19292
rect 24668 19236 24724 19246
rect 24444 19180 24668 19236
rect 24332 18452 24388 18462
rect 24332 18358 24388 18396
rect 24444 17666 24500 19180
rect 24668 19170 24724 19180
rect 25116 19236 25172 19294
rect 25116 19170 25172 19180
rect 25788 19236 25844 19246
rect 25788 19142 25844 19180
rect 24668 19010 24724 19022
rect 24668 18958 24670 19010
rect 24722 18958 24724 19010
rect 24668 18116 24724 18958
rect 25900 19012 25956 19964
rect 26572 19908 26628 21534
rect 26908 21586 26964 23996
rect 27916 24050 27972 24062
rect 27916 23998 27918 24050
rect 27970 23998 27972 24050
rect 27916 23156 27972 23998
rect 28028 24052 28084 25230
rect 37884 25284 37940 26238
rect 40236 26292 40292 26798
rect 40236 26226 40292 26236
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 25620 39956 26126
rect 39900 25554 39956 25564
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37884 25218 37940 25228
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 28364 24052 28420 24062
rect 28084 24050 28420 24052
rect 28084 23998 28366 24050
rect 28418 23998 28420 24050
rect 28084 23996 28420 23998
rect 28028 23986 28084 23996
rect 28364 23986 28420 23996
rect 27916 23090 27972 23100
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 26908 21534 26910 21586
rect 26962 21534 26964 21586
rect 26908 20914 26964 21534
rect 26908 20862 26910 20914
rect 26962 20862 26964 20914
rect 26908 20188 26964 20862
rect 26796 20132 26964 20188
rect 27020 22036 27076 22046
rect 26684 20020 26740 20030
rect 26796 20020 26852 20132
rect 26684 20018 26852 20020
rect 26684 19966 26686 20018
rect 26738 19966 26852 20018
rect 26684 19964 26852 19966
rect 26684 19954 26740 19964
rect 26348 19852 26628 19908
rect 26348 19458 26404 19852
rect 26348 19406 26350 19458
rect 26402 19406 26404 19458
rect 26348 19394 26404 19406
rect 26236 19124 26292 19134
rect 26236 19030 26292 19068
rect 26012 19012 26068 19022
rect 25900 19010 26068 19012
rect 25900 18958 26014 19010
rect 26066 18958 26068 19010
rect 25900 18956 26068 18958
rect 26012 18564 26068 18956
rect 24668 18050 24724 18060
rect 25452 18452 25508 18462
rect 24444 17614 24446 17666
rect 24498 17614 24500 17666
rect 24444 17602 24500 17614
rect 24780 17442 24836 17454
rect 24780 17390 24782 17442
rect 24834 17390 24836 17442
rect 24780 17108 24836 17390
rect 24780 17042 24836 17052
rect 24220 16930 24276 16940
rect 23772 16830 23774 16882
rect 23826 16830 23828 16882
rect 23772 16818 23828 16830
rect 23436 16718 23438 16770
rect 23490 16718 23492 16770
rect 23436 16706 23492 16718
rect 23660 16770 23716 16782
rect 23660 16718 23662 16770
rect 23714 16718 23716 16770
rect 23660 16210 23716 16718
rect 25452 16324 25508 18396
rect 26012 17666 26068 18508
rect 26012 17614 26014 17666
rect 26066 17614 26068 17666
rect 26012 17602 26068 17614
rect 26460 17668 26516 17678
rect 26460 17574 26516 17612
rect 26572 17444 26628 17454
rect 26348 17442 26628 17444
rect 26348 17390 26574 17442
rect 26626 17390 26628 17442
rect 26348 17388 26628 17390
rect 25564 17108 25620 17118
rect 26348 17108 26404 17388
rect 26572 17378 26628 17388
rect 26684 17442 26740 17454
rect 26684 17390 26686 17442
rect 26738 17390 26740 17442
rect 26684 17220 26740 17390
rect 26684 17154 26740 17164
rect 25564 17014 25620 17052
rect 25788 17052 26404 17108
rect 25788 16994 25844 17052
rect 25788 16942 25790 16994
rect 25842 16942 25844 16994
rect 25788 16930 25844 16942
rect 26796 16884 26852 19964
rect 27020 19458 27076 21980
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 27692 21474 27748 21486
rect 27692 21422 27694 21474
rect 27746 21422 27748 21474
rect 27244 20916 27300 20926
rect 27020 19406 27022 19458
rect 27074 19406 27076 19458
rect 27020 19394 27076 19406
rect 27132 20580 27188 20590
rect 27132 19458 27188 20524
rect 27132 19406 27134 19458
rect 27186 19406 27188 19458
rect 27132 19394 27188 19406
rect 27244 19460 27300 20860
rect 27692 20188 27748 21422
rect 29820 21474 29876 21486
rect 29820 21422 29822 21474
rect 29874 21422 29876 21474
rect 29484 20804 29540 20814
rect 29820 20804 29876 21422
rect 29484 20802 29876 20804
rect 29484 20750 29486 20802
rect 29538 20750 29876 20802
rect 29484 20748 29876 20750
rect 30268 21474 30324 21486
rect 30268 21422 30270 21474
rect 30322 21422 30324 21474
rect 27356 20132 27412 20142
rect 27356 20038 27412 20076
rect 27468 20132 27748 20188
rect 29148 20690 29204 20702
rect 29148 20638 29150 20690
rect 29202 20638 29204 20690
rect 27356 19460 27412 19470
rect 27244 19458 27412 19460
rect 27244 19406 27358 19458
rect 27410 19406 27412 19458
rect 27244 19404 27412 19406
rect 27356 19394 27412 19404
rect 27468 19458 27524 20132
rect 27468 19406 27470 19458
rect 27522 19406 27524 19458
rect 27468 19394 27524 19406
rect 27692 19796 27748 19806
rect 27692 18450 27748 19740
rect 29148 19796 29204 20638
rect 29260 20580 29316 20590
rect 29260 20486 29316 20524
rect 29484 20580 29540 20748
rect 29484 20514 29540 20524
rect 29148 19730 29204 19740
rect 29484 19908 29540 19918
rect 29484 19124 29540 19852
rect 29932 19908 29988 19918
rect 30268 19908 30324 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 37660 20804 37716 20814
rect 37660 20710 37716 20748
rect 29932 19906 30324 19908
rect 29932 19854 29934 19906
rect 29986 19854 30324 19906
rect 29932 19852 30324 19854
rect 29932 19842 29988 19852
rect 29484 19058 29540 19068
rect 27692 18398 27694 18450
rect 27746 18398 27748 18450
rect 27692 18386 27748 18398
rect 28028 18452 28084 18462
rect 28476 18452 28532 18462
rect 28028 18450 28532 18452
rect 28028 18398 28030 18450
rect 28082 18398 28478 18450
rect 28530 18398 28532 18450
rect 28028 18396 28532 18398
rect 28028 18386 28084 18396
rect 28476 18386 28532 18396
rect 28700 18452 28756 18462
rect 28700 18358 28756 18396
rect 29820 18452 29876 18462
rect 27692 18226 27748 18238
rect 27692 18174 27694 18226
rect 27746 18174 27748 18226
rect 27692 16994 27748 18174
rect 28364 18226 28420 18238
rect 28364 18174 28366 18226
rect 28418 18174 28420 18226
rect 27692 16942 27694 16994
rect 27746 16942 27748 16994
rect 27692 16930 27748 16942
rect 28140 17668 28196 17678
rect 27020 16884 27076 16894
rect 26796 16882 27188 16884
rect 26796 16830 27022 16882
rect 27074 16830 27188 16882
rect 26796 16828 27188 16830
rect 27020 16818 27076 16828
rect 25676 16772 25732 16782
rect 25676 16770 26068 16772
rect 25676 16718 25678 16770
rect 25730 16718 26068 16770
rect 25676 16716 26068 16718
rect 25676 16706 25732 16716
rect 25452 16268 25844 16324
rect 23660 16158 23662 16210
rect 23714 16158 23716 16210
rect 23660 16146 23716 16158
rect 25788 16212 25844 16268
rect 25788 16118 25844 16156
rect 22988 16098 23044 16110
rect 22988 16046 22990 16098
rect 23042 16046 23044 16098
rect 22988 15316 23044 16046
rect 26012 15426 26068 16716
rect 26572 16212 26628 16222
rect 26572 16100 26628 16156
rect 26572 16098 26852 16100
rect 26572 16046 26574 16098
rect 26626 16046 26852 16098
rect 26572 16044 26852 16046
rect 26572 16034 26628 16044
rect 26012 15374 26014 15426
rect 26066 15374 26068 15426
rect 26012 15362 26068 15374
rect 26348 15874 26404 15886
rect 26348 15822 26350 15874
rect 26402 15822 26404 15874
rect 23324 15316 23380 15326
rect 22988 15260 23324 15316
rect 23324 15222 23380 15260
rect 25340 15316 25396 15326
rect 25340 15222 25396 15260
rect 22876 15204 22932 15214
rect 22540 15202 22932 15204
rect 22540 15150 22878 15202
rect 22930 15150 22932 15202
rect 22540 15148 22932 15150
rect 22876 15138 22932 15148
rect 20748 14642 21028 14644
rect 20748 14590 20750 14642
rect 20802 14590 21028 14642
rect 20748 14588 21028 14590
rect 20748 14578 20804 14588
rect 17612 14532 17668 14542
rect 17836 14532 17892 14542
rect 17500 14530 17892 14532
rect 17500 14478 17614 14530
rect 17666 14478 17838 14530
rect 17890 14478 17892 14530
rect 17500 14476 17892 14478
rect 17612 14466 17668 14476
rect 17836 14466 17892 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 26348 8428 26404 15822
rect 26796 15204 26852 16044
rect 27132 15874 27188 16828
rect 27132 15822 27134 15874
rect 27186 15822 27188 15874
rect 27132 15316 27188 15822
rect 27132 15250 27188 15260
rect 26796 15148 26964 15204
rect 16828 8372 17108 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17052 3554 17108 8372
rect 25788 8372 26404 8428
rect 26908 8428 26964 15148
rect 28140 15202 28196 17612
rect 28364 17220 28420 18174
rect 28364 17154 28420 17164
rect 29820 16884 29876 18396
rect 30268 16884 30324 19852
rect 37884 19908 37940 21534
rect 39900 21474 39956 21486
rect 39900 21422 39902 21474
rect 39954 21422 39956 21474
rect 39900 20916 39956 21422
rect 39900 20850 39956 20860
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 37884 19842 37940 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37884 18450 37940 18462
rect 37884 18398 37886 18450
rect 37938 18398 37940 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 29820 16770 29876 16828
rect 29820 16718 29822 16770
rect 29874 16718 29876 16770
rect 29820 16706 29876 16718
rect 30156 16882 30324 16884
rect 30156 16830 30270 16882
rect 30322 16830 30324 16882
rect 30156 16828 30324 16830
rect 28588 15316 28644 15326
rect 28588 15222 28644 15260
rect 30044 15316 30100 15326
rect 30156 15316 30212 16828
rect 30268 16818 30324 16828
rect 37884 16884 37940 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37884 16818 37940 16828
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 40012 16884 40068 17726
rect 40012 16818 40068 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 30100 15260 30212 15316
rect 30044 15250 30100 15260
rect 28140 15150 28142 15202
rect 28194 15150 28196 15202
rect 28140 15138 28196 15150
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 26908 8372 27188 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 25788 4338 25844 8372
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 25564 4116 25620 4126
rect 17052 3502 17054 3554
rect 17106 3502 17108 3554
rect 17052 3490 17108 3502
rect 23548 3668 23604 3678
rect 16828 3444 16884 3454
rect 16828 800 16884 3388
rect 18060 3444 18116 3454
rect 18060 3330 18116 3388
rect 18060 3278 18062 3330
rect 18114 3278 18116 3330
rect 18060 3266 18116 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 23548 800 23604 3612
rect 24780 3668 24836 3678
rect 24780 3574 24836 3612
rect 25564 800 25620 4060
rect 26796 4116 26852 4126
rect 26796 4022 26852 4060
rect 27132 3554 27188 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 27132 3502 27134 3554
rect 27186 3502 27188 3554
rect 27132 3490 27188 3502
rect 16800 0 16912 800
rect 23520 0 23632 800
rect 25536 0 25648 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 16828 38220 16884 38276
rect 18060 38274 18116 38276
rect 18060 38222 18062 38274
rect 18062 38222 18114 38274
rect 18114 38222 18116 38274
rect 18060 38220 18116 38222
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4172 26908 4228 26964
rect 1932 24892 1988 24948
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1932 23548 1988 23604
rect 13132 26178 13188 26180
rect 13132 26126 13134 26178
rect 13134 26126 13186 26178
rect 13186 26126 13188 26178
rect 13132 26124 13188 26126
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 9996 25618 10052 25620
rect 9996 25566 9998 25618
rect 9998 25566 10050 25618
rect 10050 25566 10052 25618
rect 9996 25564 10052 25566
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 16716 26236 16772 26292
rect 13916 26124 13972 26180
rect 13804 25676 13860 25732
rect 12124 25394 12180 25396
rect 12124 25342 12126 25394
rect 12126 25342 12178 25394
rect 12178 25342 12180 25394
rect 12124 25340 12180 25342
rect 12684 25228 12740 25284
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 10892 24610 10948 24612
rect 10892 24558 10894 24610
rect 10894 24558 10946 24610
rect 10946 24558 10948 24610
rect 10892 24556 10948 24558
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 10892 24108 10948 24164
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 13692 25228 13748 25284
rect 14252 25564 14308 25620
rect 14028 25394 14084 25396
rect 14028 25342 14030 25394
rect 14030 25342 14082 25394
rect 14082 25342 14084 25394
rect 14028 25340 14084 25342
rect 21532 38220 21588 38276
rect 22428 38274 22484 38276
rect 22428 38222 22430 38274
rect 22430 38222 22482 38274
rect 22482 38222 22484 38274
rect 22428 38220 22484 38222
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 24220 38220 24276 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19516 37436 19572 37492
rect 20748 37490 20804 37492
rect 20748 37438 20750 37490
rect 20750 37438 20802 37490
rect 20802 37438 20804 37490
rect 20748 37436 20804 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18956 26796 19012 26852
rect 17276 26236 17332 26292
rect 16940 26124 16996 26180
rect 15148 25228 15204 25284
rect 13916 24556 13972 24612
rect 14812 24610 14868 24612
rect 14812 24558 14814 24610
rect 14814 24558 14866 24610
rect 14866 24558 14868 24610
rect 14812 24556 14868 24558
rect 14252 24444 14308 24500
rect 13692 23884 13748 23940
rect 12908 23324 12964 23380
rect 14140 24108 14196 24164
rect 13916 23378 13972 23380
rect 13916 23326 13918 23378
rect 13918 23326 13970 23378
rect 13970 23326 13972 23378
rect 13916 23324 13972 23326
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 12908 21756 12964 21812
rect 9996 21644 10052 21700
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 4172 21420 4228 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 9996 21084 10052 21140
rect 1932 20860 1988 20916
rect 12124 20860 12180 20916
rect 4284 20802 4340 20804
rect 4284 20750 4286 20802
rect 4286 20750 4338 20802
rect 4338 20750 4340 20802
rect 4284 20748 4340 20750
rect 2044 20188 2100 20244
rect 16268 25282 16324 25284
rect 16268 25230 16270 25282
rect 16270 25230 16322 25282
rect 16322 25230 16324 25282
rect 16268 25228 16324 25230
rect 16828 25228 16884 25284
rect 16156 24108 16212 24164
rect 15484 23324 15540 23380
rect 15708 23266 15764 23268
rect 15708 23214 15710 23266
rect 15710 23214 15762 23266
rect 15762 23214 15764 23266
rect 15708 23212 15764 23214
rect 17500 26178 17556 26180
rect 17500 26126 17502 26178
rect 17502 26126 17554 26178
rect 17554 26126 17556 26178
rect 17500 26124 17556 26126
rect 17948 25340 18004 25396
rect 16940 24556 16996 24612
rect 14364 21868 14420 21924
rect 16044 23884 16100 23940
rect 14140 21810 14196 21812
rect 14140 21758 14142 21810
rect 14142 21758 14194 21810
rect 14194 21758 14196 21810
rect 14140 21756 14196 21758
rect 15036 21756 15092 21812
rect 13468 21308 13524 21364
rect 13580 21532 13636 21588
rect 13244 21084 13300 21140
rect 13356 20860 13412 20916
rect 14924 21586 14980 21588
rect 14924 21534 14926 21586
rect 14926 21534 14978 21586
rect 14978 21534 14980 21586
rect 14924 21532 14980 21534
rect 14364 21308 14420 21364
rect 12572 20130 12628 20132
rect 12572 20078 12574 20130
rect 12574 20078 12626 20130
rect 12626 20078 12628 20130
rect 12572 20076 12628 20078
rect 4284 20018 4340 20020
rect 4284 19966 4286 20018
rect 4286 19966 4338 20018
rect 4338 19966 4340 20018
rect 4284 19964 4340 19966
rect 13020 19964 13076 20020
rect 1932 19794 1988 19796
rect 1932 19742 1934 19794
rect 1934 19742 1986 19794
rect 1986 19742 1988 19794
rect 1932 19740 1988 19742
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 14028 20690 14084 20692
rect 14028 20638 14030 20690
rect 14030 20638 14082 20690
rect 14082 20638 14084 20690
rect 14028 20636 14084 20638
rect 15148 21698 15204 21700
rect 15148 21646 15150 21698
rect 15150 21646 15202 21698
rect 15202 21646 15204 21698
rect 15148 21644 15204 21646
rect 15260 21308 15316 21364
rect 15148 20914 15204 20916
rect 15148 20862 15150 20914
rect 15150 20862 15202 20914
rect 15202 20862 15204 20914
rect 15148 20860 15204 20862
rect 13804 19628 13860 19684
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 10332 17612 10388 17668
rect 1932 16828 1988 16884
rect 12572 17666 12628 17668
rect 12572 17614 12574 17666
rect 12574 17614 12626 17666
rect 12626 17614 12628 17666
rect 12572 17612 12628 17614
rect 12796 17554 12852 17556
rect 12796 17502 12798 17554
rect 12798 17502 12850 17554
rect 12850 17502 12852 17554
rect 12796 17500 12852 17502
rect 12460 17388 12516 17444
rect 13356 17666 13412 17668
rect 13356 17614 13358 17666
rect 13358 17614 13410 17666
rect 13410 17614 13412 17666
rect 13356 17612 13412 17614
rect 14476 18396 14532 18452
rect 16828 23772 16884 23828
rect 15932 21868 15988 21924
rect 15708 20914 15764 20916
rect 15708 20862 15710 20914
rect 15710 20862 15762 20914
rect 15762 20862 15764 20914
rect 15708 20860 15764 20862
rect 16492 20076 16548 20132
rect 15596 19740 15652 19796
rect 13244 16882 13300 16884
rect 13244 16830 13246 16882
rect 13246 16830 13298 16882
rect 13298 16830 13300 16882
rect 13244 16828 13300 16830
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4284 16268 4340 16324
rect 1932 16156 1988 16212
rect 13580 17442 13636 17444
rect 13580 17390 13582 17442
rect 13582 17390 13634 17442
rect 13634 17390 13636 17442
rect 13580 17388 13636 17390
rect 13356 16156 13412 16212
rect 9996 16044 10052 16100
rect 12124 15986 12180 15988
rect 12124 15934 12126 15986
rect 12126 15934 12178 15986
rect 12178 15934 12180 15986
rect 12124 15932 12180 15934
rect 13692 16828 13748 16884
rect 14700 18172 14756 18228
rect 14812 18060 14868 18116
rect 16268 20018 16324 20020
rect 16268 19966 16270 20018
rect 16270 19966 16322 20018
rect 16322 19966 16324 20018
rect 16268 19964 16324 19966
rect 16268 19794 16324 19796
rect 16268 19742 16270 19794
rect 16270 19742 16322 19794
rect 16322 19742 16324 19794
rect 16268 19740 16324 19742
rect 18508 26290 18564 26292
rect 18508 26238 18510 26290
rect 18510 26238 18562 26290
rect 18562 26238 18564 26290
rect 18508 26236 18564 26238
rect 19292 26236 19348 26292
rect 18620 26124 18676 26180
rect 19180 25676 19236 25732
rect 18284 23548 18340 23604
rect 17388 23378 17444 23380
rect 17388 23326 17390 23378
rect 17390 23326 17442 23378
rect 17442 23326 17444 23378
rect 17388 23324 17444 23326
rect 18284 23266 18340 23268
rect 18284 23214 18286 23266
rect 18286 23214 18338 23266
rect 18338 23214 18340 23266
rect 18284 23212 18340 23214
rect 18508 25340 18564 25396
rect 16604 19906 16660 19908
rect 16604 19854 16606 19906
rect 16606 19854 16658 19906
rect 16658 19854 16660 19906
rect 16604 19852 16660 19854
rect 16492 19740 16548 19796
rect 17276 22370 17332 22372
rect 17276 22318 17278 22370
rect 17278 22318 17330 22370
rect 17330 22318 17332 22370
rect 17276 22316 17332 22318
rect 17612 22316 17668 22372
rect 17948 22370 18004 22372
rect 17948 22318 17950 22370
rect 17950 22318 18002 22370
rect 18002 22318 18004 22370
rect 17948 22316 18004 22318
rect 18284 22204 18340 22260
rect 17948 21868 18004 21924
rect 17500 21474 17556 21476
rect 17500 21422 17502 21474
rect 17502 21422 17554 21474
rect 17554 21422 17556 21474
rect 17500 21420 17556 21422
rect 18060 21474 18116 21476
rect 18060 21422 18062 21474
rect 18062 21422 18114 21474
rect 18114 21422 18116 21474
rect 18060 21420 18116 21422
rect 18060 21196 18116 21252
rect 16828 19068 16884 19124
rect 16380 18956 16436 19012
rect 15820 18396 15876 18452
rect 15036 18284 15092 18340
rect 14028 16882 14084 16884
rect 14028 16830 14030 16882
rect 14030 16830 14082 16882
rect 14082 16830 14084 16882
rect 14028 16828 14084 16830
rect 13804 16098 13860 16100
rect 13804 16046 13806 16098
rect 13806 16046 13858 16098
rect 13858 16046 13860 16098
rect 13804 16044 13860 16046
rect 14028 16098 14084 16100
rect 14028 16046 14030 16098
rect 14030 16046 14082 16098
rect 14082 16046 14084 16098
rect 14028 16044 14084 16046
rect 16156 18284 16212 18340
rect 16044 18226 16100 18228
rect 16044 18174 16046 18226
rect 16046 18174 16098 18226
rect 16098 18174 16100 18226
rect 16044 18172 16100 18174
rect 16156 17836 16212 17892
rect 16828 17500 16884 17556
rect 16940 16156 16996 16212
rect 16380 16098 16436 16100
rect 16380 16046 16382 16098
rect 16382 16046 16434 16098
rect 16434 16046 16436 16098
rect 16380 16044 16436 16046
rect 17052 18396 17108 18452
rect 19068 25228 19124 25284
rect 18956 23772 19012 23828
rect 19852 26962 19908 26964
rect 19852 26910 19854 26962
rect 19854 26910 19906 26962
rect 19906 26910 19908 26962
rect 19852 26908 19908 26910
rect 20300 26908 20356 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20076 25676 20132 25732
rect 19292 25340 19348 25396
rect 20188 25340 20244 25396
rect 19516 24668 19572 24724
rect 19740 25282 19796 25284
rect 19740 25230 19742 25282
rect 19742 25230 19794 25282
rect 19794 25230 19796 25282
rect 19740 25228 19796 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19852 24946 19908 24948
rect 19852 24894 19854 24946
rect 19854 24894 19906 24946
rect 19906 24894 19908 24946
rect 19852 24892 19908 24894
rect 20748 26850 20804 26852
rect 20748 26798 20750 26850
rect 20750 26798 20802 26850
rect 20802 26798 20804 26850
rect 20748 26796 20804 26798
rect 21532 27074 21588 27076
rect 21532 27022 21534 27074
rect 21534 27022 21586 27074
rect 21586 27022 21588 27074
rect 21532 27020 21588 27022
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 40236 36370 40292 36372
rect 40236 36318 40238 36370
rect 40238 36318 40290 36370
rect 40290 36318 40292 36370
rect 40236 36316 40292 36318
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 24108 27020 24164 27076
rect 22204 26684 22260 26740
rect 21532 25228 21588 25284
rect 22876 26290 22932 26292
rect 22876 26238 22878 26290
rect 22878 26238 22930 26290
rect 22930 26238 22932 26290
rect 22876 26236 22932 26238
rect 22652 25228 22708 25284
rect 20300 24892 20356 24948
rect 19292 24220 19348 24276
rect 19068 23324 19124 23380
rect 19180 23660 19236 23716
rect 19292 23548 19348 23604
rect 19964 24722 20020 24724
rect 19964 24670 19966 24722
rect 19966 24670 20018 24722
rect 20018 24670 20020 24722
rect 19964 24668 20020 24670
rect 21308 24668 21364 24724
rect 19740 24220 19796 24276
rect 19516 23772 19572 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19292 22316 19348 22372
rect 19068 21810 19124 21812
rect 19068 21758 19070 21810
rect 19070 21758 19122 21810
rect 19122 21758 19124 21810
rect 19068 21756 19124 21758
rect 19404 21586 19460 21588
rect 19404 21534 19406 21586
rect 19406 21534 19458 21586
rect 19458 21534 19460 21586
rect 19404 21532 19460 21534
rect 18844 21420 18900 21476
rect 18620 20636 18676 20692
rect 19404 20636 19460 20692
rect 18396 19852 18452 19908
rect 17724 19122 17780 19124
rect 17724 19070 17726 19122
rect 17726 19070 17778 19122
rect 17778 19070 17780 19122
rect 17724 19068 17780 19070
rect 17836 19010 17892 19012
rect 17836 18958 17838 19010
rect 17838 18958 17890 19010
rect 17890 18958 17892 19010
rect 17836 18956 17892 18958
rect 17276 18396 17332 18452
rect 14476 15986 14532 15988
rect 14476 15934 14478 15986
rect 14478 15934 14530 15986
rect 14530 15934 14532 15986
rect 14476 15932 14532 15934
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 17612 18060 17668 18116
rect 17724 17612 17780 17668
rect 18508 19964 18564 20020
rect 18844 19794 18900 19796
rect 18844 19742 18846 19794
rect 18846 19742 18898 19794
rect 18898 19742 18900 19794
rect 18844 19740 18900 19742
rect 19516 20076 19572 20132
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20188 21756 20244 21812
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19628 19794 19684 19796
rect 19628 19742 19630 19794
rect 19630 19742 19682 19794
rect 19682 19742 19684 19794
rect 19628 19740 19684 19742
rect 19516 19180 19572 19236
rect 20636 23548 20692 23604
rect 20412 22092 20468 22148
rect 21532 23548 21588 23604
rect 21308 22258 21364 22260
rect 21308 22206 21310 22258
rect 21310 22206 21362 22258
rect 21362 22206 21364 22258
rect 21308 22204 21364 22206
rect 20748 21756 20804 21812
rect 21196 21756 21252 21812
rect 20300 19964 20356 20020
rect 20412 21420 20468 21476
rect 20188 19180 20244 19236
rect 20524 20300 20580 20356
rect 19964 18956 20020 19012
rect 18284 17948 18340 18004
rect 18060 17890 18116 17892
rect 18060 17838 18062 17890
rect 18062 17838 18114 17890
rect 18114 17838 18116 17890
rect 18060 17836 18116 17838
rect 19068 18450 19124 18452
rect 19068 18398 19070 18450
rect 19070 18398 19122 18450
rect 19122 18398 19124 18450
rect 19068 18396 19124 18398
rect 19068 18060 19124 18116
rect 17388 17554 17444 17556
rect 17388 17502 17390 17554
rect 17390 17502 17442 17554
rect 17442 17502 17444 17554
rect 17388 17500 17444 17502
rect 18732 17554 18788 17556
rect 18732 17502 18734 17554
rect 18734 17502 18786 17554
rect 18786 17502 18788 17554
rect 18732 17500 18788 17502
rect 19404 17836 19460 17892
rect 20860 20130 20916 20132
rect 20860 20078 20862 20130
rect 20862 20078 20914 20130
rect 20914 20078 20916 20130
rect 20860 20076 20916 20078
rect 20748 19234 20804 19236
rect 20748 19182 20750 19234
rect 20750 19182 20802 19234
rect 20802 19182 20804 19234
rect 20748 19180 20804 19182
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20972 19180 21028 19236
rect 19852 18338 19908 18340
rect 19852 18286 19854 18338
rect 19854 18286 19906 18338
rect 19906 18286 19908 18338
rect 19852 18284 19908 18286
rect 20188 18172 20244 18228
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20636 17890 20692 17892
rect 20636 17838 20638 17890
rect 20638 17838 20690 17890
rect 20690 17838 20692 17890
rect 20636 17836 20692 17838
rect 20748 17554 20804 17556
rect 20748 17502 20750 17554
rect 20750 17502 20802 17554
rect 20802 17502 20804 17554
rect 20748 17500 20804 17502
rect 19852 17052 19908 17108
rect 18396 16940 18452 16996
rect 17948 16882 18004 16884
rect 17948 16830 17950 16882
rect 17950 16830 18002 16882
rect 18002 16830 18004 16882
rect 17948 16828 18004 16830
rect 19404 16940 19460 16996
rect 19180 16882 19236 16884
rect 19180 16830 19182 16882
rect 19182 16830 19234 16882
rect 19234 16830 19236 16882
rect 19180 16828 19236 16830
rect 18508 16716 18564 16772
rect 20076 16828 20132 16884
rect 19964 16716 20020 16772
rect 18508 16044 18564 16100
rect 14700 14700 14756 14756
rect 15708 14754 15764 14756
rect 15708 14702 15710 14754
rect 15710 14702 15762 14754
rect 15762 14702 15764 14754
rect 15708 14700 15764 14702
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20076 15314 20132 15316
rect 20076 15262 20078 15314
rect 20078 15262 20130 15314
rect 20130 15262 20132 15314
rect 20076 15260 20132 15262
rect 21308 20300 21364 20356
rect 21308 20076 21364 20132
rect 22764 23772 22820 23828
rect 23324 25228 23380 25284
rect 24780 27074 24836 27076
rect 24780 27022 24782 27074
rect 24782 27022 24834 27074
rect 24834 27022 24836 27074
rect 24780 27020 24836 27022
rect 24332 26236 24388 26292
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 23212 23714 23268 23716
rect 23212 23662 23214 23714
rect 23214 23662 23266 23714
rect 23266 23662 23268 23714
rect 23212 23660 23268 23662
rect 26908 25618 26964 25620
rect 26908 25566 26910 25618
rect 26910 25566 26962 25618
rect 26962 25566 26964 25618
rect 26908 25564 26964 25566
rect 24108 24108 24164 24164
rect 25340 25228 25396 25284
rect 24668 24444 24724 24500
rect 25004 24108 25060 24164
rect 23996 23660 24052 23716
rect 23100 23436 23156 23492
rect 22204 23100 22260 23156
rect 22092 22204 22148 22260
rect 22316 21756 22372 21812
rect 21980 20914 22036 20916
rect 21980 20862 21982 20914
rect 21982 20862 22034 20914
rect 22034 20862 22036 20914
rect 21980 20860 22036 20862
rect 23324 23154 23380 23156
rect 23324 23102 23326 23154
rect 23326 23102 23378 23154
rect 23378 23102 23380 23154
rect 23324 23100 23380 23102
rect 22876 21868 22932 21924
rect 23100 21644 23156 21700
rect 23324 20802 23380 20804
rect 23324 20750 23326 20802
rect 23326 20750 23378 20802
rect 23378 20750 23380 20802
rect 23324 20748 23380 20750
rect 22428 20076 22484 20132
rect 21868 19964 21924 20020
rect 21308 19180 21364 19236
rect 22540 20018 22596 20020
rect 22540 19966 22542 20018
rect 22542 19966 22594 20018
rect 22594 19966 22596 20018
rect 22540 19964 22596 19966
rect 23772 20018 23828 20020
rect 23772 19966 23774 20018
rect 23774 19966 23826 20018
rect 23826 19966 23828 20018
rect 23772 19964 23828 19966
rect 22764 19852 22820 19908
rect 23548 19906 23604 19908
rect 23548 19854 23550 19906
rect 23550 19854 23602 19906
rect 23602 19854 23604 19906
rect 23548 19852 23604 19854
rect 21308 18956 21364 19012
rect 21532 18450 21588 18452
rect 21532 18398 21534 18450
rect 21534 18398 21586 18450
rect 21586 18398 21588 18450
rect 21532 18396 21588 18398
rect 21084 16994 21140 16996
rect 21084 16942 21086 16994
rect 21086 16942 21138 16994
rect 21138 16942 21140 16994
rect 21084 16940 21140 16942
rect 21980 19068 22036 19124
rect 22316 18450 22372 18452
rect 22316 18398 22318 18450
rect 22318 18398 22370 18450
rect 22370 18398 22372 18450
rect 22316 18396 22372 18398
rect 22204 18060 22260 18116
rect 23212 18508 23268 18564
rect 22764 18172 22820 18228
rect 22988 18396 23044 18452
rect 22988 17666 23044 17668
rect 22988 17614 22990 17666
rect 22990 17614 23042 17666
rect 23042 17614 23044 17666
rect 22988 17612 23044 17614
rect 22540 17500 22596 17556
rect 23884 18562 23940 18564
rect 23884 18510 23886 18562
rect 23886 18510 23938 18562
rect 23938 18510 23940 18562
rect 23884 18508 23940 18510
rect 23772 18396 23828 18452
rect 23324 18284 23380 18340
rect 23772 18172 23828 18228
rect 24108 19794 24164 19796
rect 24108 19742 24110 19794
rect 24110 19742 24162 19794
rect 24162 19742 24164 19794
rect 24108 19740 24164 19742
rect 24108 18060 24164 18116
rect 23996 17948 24052 18004
rect 23772 17052 23828 17108
rect 25004 23660 25060 23716
rect 24444 22092 24500 22148
rect 24332 21868 24388 21924
rect 24444 21756 24500 21812
rect 24780 21532 24836 21588
rect 25004 22146 25060 22148
rect 25004 22094 25006 22146
rect 25006 22094 25058 22146
rect 25058 22094 25060 22146
rect 25004 22092 25060 22094
rect 25228 22092 25284 22148
rect 25564 24834 25620 24836
rect 25564 24782 25566 24834
rect 25566 24782 25618 24834
rect 25618 24782 25620 24834
rect 25564 24780 25620 24782
rect 27356 25564 27412 25620
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 27580 25282 27636 25284
rect 27580 25230 27582 25282
rect 27582 25230 27634 25282
rect 27634 25230 27636 25282
rect 27580 25228 27636 25230
rect 26908 24780 26964 24836
rect 25452 24498 25508 24500
rect 25452 24446 25454 24498
rect 25454 24446 25506 24498
rect 25506 24446 25508 24498
rect 25452 24444 25508 24446
rect 26908 23996 26964 24052
rect 25452 23436 25508 23492
rect 26124 23100 26180 23156
rect 25676 22258 25732 22260
rect 25676 22206 25678 22258
rect 25678 22206 25730 22258
rect 25730 22206 25732 22258
rect 25676 22204 25732 22206
rect 25900 21868 25956 21924
rect 25564 21810 25620 21812
rect 25564 21758 25566 21810
rect 25566 21758 25618 21810
rect 25618 21758 25620 21810
rect 25564 21756 25620 21758
rect 25452 21644 25508 21700
rect 26236 21586 26292 21588
rect 26236 21534 26238 21586
rect 26238 21534 26290 21586
rect 26290 21534 26292 21586
rect 26236 21532 26292 21534
rect 26012 20860 26068 20916
rect 26460 20076 26516 20132
rect 24668 19180 24724 19236
rect 24332 18450 24388 18452
rect 24332 18398 24334 18450
rect 24334 18398 24386 18450
rect 24386 18398 24388 18450
rect 24332 18396 24388 18398
rect 25116 19180 25172 19236
rect 25788 19234 25844 19236
rect 25788 19182 25790 19234
rect 25790 19182 25842 19234
rect 25842 19182 25844 19234
rect 25788 19180 25844 19182
rect 40236 26236 40292 26292
rect 39900 25564 39956 25620
rect 37884 25228 37940 25284
rect 40012 24892 40068 24948
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 28028 23996 28084 24052
rect 27916 23100 27972 23156
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 27020 21980 27076 22036
rect 26236 19122 26292 19124
rect 26236 19070 26238 19122
rect 26238 19070 26290 19122
rect 26290 19070 26292 19122
rect 26236 19068 26292 19070
rect 26012 18508 26068 18564
rect 24668 18060 24724 18116
rect 25452 18396 25508 18452
rect 24780 17052 24836 17108
rect 24220 16940 24276 16996
rect 26460 17666 26516 17668
rect 26460 17614 26462 17666
rect 26462 17614 26514 17666
rect 26514 17614 26516 17666
rect 26460 17612 26516 17614
rect 26684 17164 26740 17220
rect 25564 17106 25620 17108
rect 25564 17054 25566 17106
rect 25566 17054 25618 17106
rect 25618 17054 25620 17106
rect 25564 17052 25620 17054
rect 27244 20860 27300 20916
rect 27132 20524 27188 20580
rect 27356 20130 27412 20132
rect 27356 20078 27358 20130
rect 27358 20078 27410 20130
rect 27410 20078 27412 20130
rect 27356 20076 27412 20078
rect 27692 19740 27748 19796
rect 29260 20578 29316 20580
rect 29260 20526 29262 20578
rect 29262 20526 29314 20578
rect 29314 20526 29316 20578
rect 29260 20524 29316 20526
rect 29484 20524 29540 20580
rect 29148 19740 29204 19796
rect 29484 19906 29540 19908
rect 29484 19854 29486 19906
rect 29486 19854 29538 19906
rect 29538 19854 29540 19906
rect 29484 19852 29540 19854
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 37660 20802 37716 20804
rect 37660 20750 37662 20802
rect 37662 20750 37714 20802
rect 37714 20750 37716 20802
rect 37660 20748 37716 20750
rect 29484 19068 29540 19124
rect 28700 18450 28756 18452
rect 28700 18398 28702 18450
rect 28702 18398 28754 18450
rect 28754 18398 28756 18450
rect 28700 18396 28756 18398
rect 29820 18396 29876 18452
rect 28140 17612 28196 17668
rect 25788 16210 25844 16212
rect 25788 16158 25790 16210
rect 25790 16158 25842 16210
rect 25842 16158 25844 16210
rect 25788 16156 25844 16158
rect 26572 16156 26628 16212
rect 23324 15314 23380 15316
rect 23324 15262 23326 15314
rect 23326 15262 23378 15314
rect 23378 15262 23380 15314
rect 23324 15260 23380 15262
rect 25340 15314 25396 15316
rect 25340 15262 25342 15314
rect 25342 15262 25394 15314
rect 25394 15262 25396 15314
rect 25340 15260 25396 15262
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 27132 15260 27188 15316
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 28364 17164 28420 17220
rect 39900 20860 39956 20916
rect 40012 20188 40068 20244
rect 37884 19852 37940 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 29820 16828 29876 16884
rect 28588 15314 28644 15316
rect 28588 15262 28590 15314
rect 28590 15262 28642 15314
rect 28642 15262 28644 15314
rect 28588 15260 28644 15262
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37884 16828 37940 16884
rect 40012 16828 40068 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 30044 15260 30100 15316
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 25564 4060 25620 4116
rect 23548 3612 23604 3668
rect 16828 3388 16884 3444
rect 18060 3388 18116 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 24780 3666 24836 3668
rect 24780 3614 24782 3666
rect 24782 3614 24834 3666
rect 24834 3614 24836 3666
rect 24780 3612 24836 3614
rect 26796 4114 26852 4116
rect 26796 4062 26798 4114
rect 26798 4062 26850 4114
rect 26850 4062 26852 4114
rect 26796 4060 26852 4062
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16818 38220 16828 38276
rect 16884 38220 18060 38276
rect 18116 38220 18126 38276
rect 21522 38220 21532 38276
rect 21588 38220 22428 38276
rect 22484 38220 22494 38276
rect 24210 38220 24220 38276
rect 24276 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 19506 37436 19516 37492
rect 19572 37436 20748 37492
rect 20804 37436 20814 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 0 36372 800 36400
rect 41200 36372 42000 36400
rect 0 36316 1708 36372
rect 1764 36316 1774 36372
rect 40226 36316 40236 36372
rect 40292 36316 42000 36372
rect 0 36288 800 36316
rect 41200 36288 42000 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 21522 27020 21532 27076
rect 21588 27020 24108 27076
rect 24164 27020 24780 27076
rect 24836 27020 24846 27076
rect 0 26964 800 26992
rect 0 26908 4172 26964
rect 4228 26908 4238 26964
rect 19842 26908 19852 26964
rect 19908 26908 20300 26964
rect 20356 26908 22260 26964
rect 0 26880 800 26908
rect 18946 26796 18956 26852
rect 19012 26796 20748 26852
rect 20804 26796 20814 26852
rect 22204 26740 22260 26908
rect 22194 26684 22204 26740
rect 22260 26684 22270 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 41200 26292 42000 26320
rect 16706 26236 16716 26292
rect 16772 26236 17276 26292
rect 17332 26236 17342 26292
rect 18498 26236 18508 26292
rect 18564 26236 19292 26292
rect 19348 26236 19358 26292
rect 22866 26236 22876 26292
rect 22932 26236 24332 26292
rect 24388 26236 24398 26292
rect 40226 26236 40236 26292
rect 40292 26236 42000 26292
rect 41200 26208 42000 26236
rect 13122 26124 13132 26180
rect 13188 26124 13916 26180
rect 13972 26124 13982 26180
rect 16930 26124 16940 26180
rect 16996 26124 17500 26180
rect 17556 26124 18620 26180
rect 18676 26124 18686 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 13794 25676 13804 25732
rect 13860 25676 19180 25732
rect 19236 25676 20076 25732
rect 20132 25676 20142 25732
rect 41200 25620 42000 25648
rect 8372 25564 9996 25620
rect 10052 25564 14252 25620
rect 14308 25564 14318 25620
rect 26898 25564 26908 25620
rect 26964 25564 27356 25620
rect 27412 25564 31948 25620
rect 39890 25564 39900 25620
rect 39956 25564 42000 25620
rect 8372 25508 8428 25564
rect 4274 25452 4284 25508
rect 4340 25452 8428 25508
rect 31892 25508 31948 25564
rect 41200 25536 42000 25564
rect 31892 25452 37660 25508
rect 37716 25452 37726 25508
rect 12114 25340 12124 25396
rect 12180 25340 14028 25396
rect 14084 25340 14094 25396
rect 17938 25340 17948 25396
rect 18004 25340 18508 25396
rect 18564 25340 19292 25396
rect 19348 25340 20188 25396
rect 20244 25340 20254 25396
rect 12674 25228 12684 25284
rect 12740 25228 13692 25284
rect 13748 25228 15148 25284
rect 15204 25228 16268 25284
rect 16324 25228 16334 25284
rect 16818 25228 16828 25284
rect 16884 25228 19068 25284
rect 19124 25228 19134 25284
rect 19730 25228 19740 25284
rect 19796 25228 21532 25284
rect 21588 25228 22652 25284
rect 22708 25228 22718 25284
rect 23314 25228 23324 25284
rect 23380 25228 25340 25284
rect 25396 25228 25406 25284
rect 27570 25228 27580 25284
rect 27636 25228 37884 25284
rect 37940 25228 37950 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 19842 24892 19852 24948
rect 19908 24892 20300 24948
rect 20356 24892 20366 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 25554 24780 25564 24836
rect 25620 24780 26908 24836
rect 26964 24780 26974 24836
rect 4274 24668 4284 24724
rect 4340 24668 8428 24724
rect 19506 24668 19516 24724
rect 19572 24668 19964 24724
rect 20020 24668 21308 24724
rect 21364 24668 21374 24724
rect 8372 24612 8428 24668
rect 8372 24556 10892 24612
rect 10948 24556 10958 24612
rect 13906 24556 13916 24612
rect 13972 24556 14812 24612
rect 14868 24556 16940 24612
rect 16996 24556 17006 24612
rect 14252 24500 14308 24556
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 14242 24444 14252 24500
rect 14308 24444 14318 24500
rect 24658 24444 24668 24500
rect 24724 24444 25452 24500
rect 25508 24444 25518 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 19282 24220 19292 24276
rect 19348 24220 19740 24276
rect 19796 24220 19806 24276
rect 0 24192 800 24220
rect 10882 24108 10892 24164
rect 10948 24108 14140 24164
rect 14196 24108 14206 24164
rect 16146 24108 16156 24164
rect 16212 24108 24108 24164
rect 24164 24108 25004 24164
rect 25060 24108 25070 24164
rect 4274 23884 4284 23940
rect 4340 23884 13692 23940
rect 13748 23884 16044 23940
rect 16100 23884 16110 23940
rect 16818 23772 16828 23828
rect 16884 23772 18956 23828
rect 19012 23772 19022 23828
rect 19506 23772 19516 23828
rect 19572 23772 22764 23828
rect 22820 23772 22830 23828
rect 26852 23716 26908 24052
rect 26964 23996 28028 24052
rect 28084 23996 28094 24052
rect 19170 23660 19180 23716
rect 19236 23660 23212 23716
rect 23268 23660 23996 23716
rect 24052 23660 25004 23716
rect 25060 23660 26908 23716
rect 0 23604 800 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 18274 23548 18284 23604
rect 18340 23548 19292 23604
rect 19348 23548 19358 23604
rect 20626 23548 20636 23604
rect 20692 23548 21532 23604
rect 21588 23548 21598 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 23090 23436 23100 23492
rect 23156 23436 25452 23492
rect 25508 23436 25518 23492
rect 23100 23380 23156 23436
rect 12898 23324 12908 23380
rect 12964 23324 13916 23380
rect 13972 23324 13982 23380
rect 15474 23324 15484 23380
rect 15540 23324 17388 23380
rect 17444 23324 17454 23380
rect 19058 23324 19068 23380
rect 19124 23324 23156 23380
rect 15698 23212 15708 23268
rect 15764 23212 18284 23268
rect 18340 23212 18350 23268
rect 22194 23100 22204 23156
rect 22260 23100 23324 23156
rect 23380 23100 23390 23156
rect 26114 23100 26124 23156
rect 26180 23100 27916 23156
rect 27972 23100 37660 23156
rect 37716 23100 37726 23156
rect 41200 22932 42000 22960
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 17266 22316 17276 22372
rect 17332 22316 17612 22372
rect 17668 22316 17948 22372
rect 18004 22316 19292 22372
rect 19348 22316 19358 22372
rect 18274 22204 18284 22260
rect 18340 22204 21308 22260
rect 21364 22204 22092 22260
rect 22148 22204 22158 22260
rect 24444 22204 25676 22260
rect 25732 22204 25742 22260
rect 24444 22148 24500 22204
rect 18060 22092 20412 22148
rect 20468 22092 24444 22148
rect 24500 22092 24510 22148
rect 24994 22092 25004 22148
rect 25060 22092 25228 22148
rect 25284 22092 26908 22148
rect 18060 22036 18116 22092
rect 26852 22036 26908 22092
rect 18050 21980 18060 22036
rect 18116 21980 18126 22036
rect 26852 21980 27020 22036
rect 27076 21980 27086 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 14354 21868 14364 21924
rect 14420 21868 15932 21924
rect 15988 21868 17948 21924
rect 18004 21868 18014 21924
rect 22866 21868 22876 21924
rect 22932 21868 24332 21924
rect 24388 21868 25900 21924
rect 25956 21868 25966 21924
rect 12898 21756 12908 21812
rect 12964 21756 14140 21812
rect 14196 21756 15036 21812
rect 15092 21756 15102 21812
rect 19058 21756 19068 21812
rect 19124 21756 20188 21812
rect 20244 21756 20748 21812
rect 20804 21756 21196 21812
rect 21252 21756 22316 21812
rect 22372 21756 22382 21812
rect 24434 21756 24444 21812
rect 24500 21756 25564 21812
rect 25620 21756 25630 21812
rect 8372 21644 9996 21700
rect 10052 21644 15148 21700
rect 15204 21644 15214 21700
rect 23090 21644 23100 21700
rect 23156 21644 25452 21700
rect 25508 21644 25518 21700
rect 8372 21588 8428 21644
rect 4274 21532 4284 21588
rect 4340 21532 8428 21588
rect 13570 21532 13580 21588
rect 13636 21532 14924 21588
rect 14980 21532 14990 21588
rect 17500 21532 19404 21588
rect 19460 21532 19470 21588
rect 24770 21532 24780 21588
rect 24836 21532 26236 21588
rect 26292 21532 26302 21588
rect 17500 21476 17556 21532
rect 4162 21420 4172 21476
rect 4228 21420 17500 21476
rect 17556 21420 17566 21476
rect 18050 21420 18060 21476
rect 18116 21420 18844 21476
rect 18900 21420 20412 21476
rect 20468 21420 20478 21476
rect 13458 21308 13468 21364
rect 13524 21308 14364 21364
rect 14420 21308 15260 21364
rect 15316 21308 15326 21364
rect 18022 21196 18060 21252
rect 18116 21196 18126 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 8372 21084 9996 21140
rect 10052 21084 13244 21140
rect 13300 21084 13310 21140
rect 0 20916 800 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 0 20832 800 20860
rect 8372 20804 8428 21084
rect 41200 20916 42000 20944
rect 12114 20860 12124 20916
rect 12180 20860 13356 20916
rect 13412 20860 13422 20916
rect 15138 20860 15148 20916
rect 15204 20860 15708 20916
rect 15764 20860 15774 20916
rect 21970 20860 21980 20916
rect 22036 20860 26012 20916
rect 26068 20860 27244 20916
rect 27300 20860 27310 20916
rect 39890 20860 39900 20916
rect 39956 20860 42000 20916
rect 41200 20832 42000 20860
rect 4274 20748 4284 20804
rect 4340 20748 8428 20804
rect 20066 20748 20076 20804
rect 20132 20748 23324 20804
rect 23380 20748 23390 20804
rect 31892 20748 37660 20804
rect 37716 20748 37726 20804
rect 14018 20636 14028 20692
rect 14084 20636 18620 20692
rect 18676 20636 19404 20692
rect 19460 20636 19470 20692
rect 31892 20580 31948 20748
rect 27122 20524 27132 20580
rect 27188 20524 29260 20580
rect 29316 20524 29326 20580
rect 29474 20524 29484 20580
rect 29540 20524 31948 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 20514 20300 20524 20356
rect 20580 20300 21308 20356
rect 21364 20300 21374 20356
rect 0 20244 800 20272
rect 41200 20244 42000 20272
rect 0 20188 2044 20244
rect 2100 20188 2110 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 0 20160 800 20188
rect 41200 20160 42000 20188
rect 12562 20076 12572 20132
rect 12628 20076 16492 20132
rect 16548 20076 16558 20132
rect 19506 20076 19516 20132
rect 19572 20076 20860 20132
rect 20916 20076 20926 20132
rect 21298 20076 21308 20132
rect 21364 20076 22428 20132
rect 22484 20076 22494 20132
rect 26450 20076 26460 20132
rect 26516 20076 27356 20132
rect 27412 20076 27422 20132
rect 4274 19964 4284 20020
rect 4340 19964 13020 20020
rect 13076 19964 16268 20020
rect 16324 19964 16334 20020
rect 18498 19964 18508 20020
rect 18564 19964 20300 20020
rect 20356 19964 20366 20020
rect 21858 19964 21868 20020
rect 21924 19964 22540 20020
rect 22596 19964 23772 20020
rect 23828 19964 23838 20020
rect 20300 19908 20356 19964
rect 16594 19852 16604 19908
rect 16660 19852 18396 19908
rect 18452 19852 18462 19908
rect 20300 19852 22764 19908
rect 22820 19852 23548 19908
rect 23604 19852 23614 19908
rect 29474 19852 29484 19908
rect 29540 19852 37884 19908
rect 37940 19852 37950 19908
rect 1922 19740 1932 19796
rect 1988 19740 1998 19796
rect 15586 19740 15596 19796
rect 15652 19740 16268 19796
rect 16324 19740 16334 19796
rect 16482 19740 16492 19796
rect 16548 19740 18844 19796
rect 18900 19740 18910 19796
rect 19618 19740 19628 19796
rect 19684 19740 19694 19796
rect 24098 19740 24108 19796
rect 24164 19740 27692 19796
rect 27748 19740 29148 19796
rect 29204 19740 29214 19796
rect 0 19572 800 19600
rect 1932 19572 1988 19740
rect 19628 19684 19684 19740
rect 13794 19628 13804 19684
rect 13860 19628 19684 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 0 19516 1988 19572
rect 0 19488 800 19516
rect 19506 19180 19516 19236
rect 19572 19180 20188 19236
rect 20244 19180 20254 19236
rect 20738 19180 20748 19236
rect 20804 19180 20972 19236
rect 21028 19180 21308 19236
rect 21364 19180 21374 19236
rect 24658 19180 24668 19236
rect 24724 19180 25116 19236
rect 25172 19180 25788 19236
rect 25844 19180 25854 19236
rect 16818 19068 16828 19124
rect 16884 19068 17724 19124
rect 17780 19068 21980 19124
rect 22036 19068 22046 19124
rect 26226 19068 26236 19124
rect 26292 19068 29484 19124
rect 29540 19068 29550 19124
rect 16370 18956 16380 19012
rect 16436 18956 17836 19012
rect 17892 18956 17902 19012
rect 19954 18956 19964 19012
rect 20020 18956 21308 19012
rect 21364 18956 21374 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 23202 18508 23212 18564
rect 23268 18508 23884 18564
rect 23940 18508 26012 18564
rect 26068 18508 26078 18564
rect 14466 18396 14476 18452
rect 14532 18396 15820 18452
rect 15876 18396 17052 18452
rect 17108 18396 17118 18452
rect 17266 18396 17276 18452
rect 17332 18396 19068 18452
rect 19124 18396 19134 18452
rect 21522 18396 21532 18452
rect 21588 18396 22316 18452
rect 22372 18396 22382 18452
rect 22978 18396 22988 18452
rect 23044 18396 23772 18452
rect 23828 18396 23838 18452
rect 24322 18396 24332 18452
rect 24388 18396 25452 18452
rect 25508 18396 25518 18452
rect 28690 18396 28700 18452
rect 28756 18396 29820 18452
rect 29876 18396 29886 18452
rect 15026 18284 15036 18340
rect 15092 18284 16156 18340
rect 16212 18284 16222 18340
rect 19842 18284 19852 18340
rect 19908 18284 23324 18340
rect 23380 18284 23390 18340
rect 41200 18228 42000 18256
rect 14690 18172 14700 18228
rect 14756 18172 16044 18228
rect 16100 18172 16110 18228
rect 20178 18172 20188 18228
rect 20244 18172 22764 18228
rect 22820 18172 23772 18228
rect 23828 18172 23838 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 14802 18060 14812 18116
rect 14868 18060 17612 18116
rect 17668 18060 17678 18116
rect 19058 18060 19068 18116
rect 19124 18060 22204 18116
rect 22260 18060 24108 18116
rect 24164 18060 24668 18116
rect 24724 18060 24734 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 18274 17948 18284 18004
rect 18340 17948 23996 18004
rect 24052 17948 24062 18004
rect 16146 17836 16156 17892
rect 16212 17836 18060 17892
rect 18116 17836 18126 17892
rect 19394 17836 19404 17892
rect 19460 17836 20636 17892
rect 20692 17836 20702 17892
rect 4274 17612 4284 17668
rect 4340 17612 10332 17668
rect 10388 17612 10398 17668
rect 12562 17612 12572 17668
rect 12628 17612 13356 17668
rect 13412 17612 13422 17668
rect 17714 17612 17724 17668
rect 17780 17612 22988 17668
rect 23044 17612 23054 17668
rect 26450 17612 26460 17668
rect 26516 17612 28140 17668
rect 28196 17612 37660 17668
rect 37716 17612 37726 17668
rect 10332 17556 10388 17612
rect 10332 17500 12796 17556
rect 12852 17500 12862 17556
rect 16818 17500 16828 17556
rect 16884 17500 17388 17556
rect 17444 17500 18732 17556
rect 18788 17500 18798 17556
rect 20738 17500 20748 17556
rect 20804 17500 22540 17556
rect 22596 17500 22606 17556
rect 12450 17388 12460 17444
rect 12516 17388 13580 17444
rect 13636 17388 13646 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 20188 17164 26684 17220
rect 26740 17164 28364 17220
rect 28420 17164 28430 17220
rect 20188 17108 20244 17164
rect 19842 17052 19852 17108
rect 19908 17052 20244 17108
rect 23762 17052 23772 17108
rect 23828 17052 24780 17108
rect 24836 17052 25564 17108
rect 25620 17052 25630 17108
rect 18386 16940 18396 16996
rect 18452 16940 19404 16996
rect 19460 16940 21084 16996
rect 21140 16940 24220 16996
rect 24276 16940 24286 16996
rect 0 16884 800 16912
rect 41200 16884 42000 16912
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 13234 16828 13244 16884
rect 13300 16828 13692 16884
rect 13748 16828 14028 16884
rect 14084 16828 14094 16884
rect 17938 16828 17948 16884
rect 18004 16828 19180 16884
rect 19236 16828 20076 16884
rect 20132 16828 20142 16884
rect 29810 16828 29820 16884
rect 29876 16828 37884 16884
rect 37940 16828 37950 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 0 16800 800 16828
rect 41200 16800 42000 16828
rect 18498 16716 18508 16772
rect 18564 16716 19964 16772
rect 20020 16716 20030 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 4274 16268 4284 16324
rect 4340 16268 8428 16324
rect 0 16212 800 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 0 16128 800 16156
rect 8372 16100 8428 16268
rect 13346 16156 13356 16212
rect 13412 16156 16940 16212
rect 16996 16156 17006 16212
rect 25778 16156 25788 16212
rect 25844 16156 26572 16212
rect 26628 16156 26638 16212
rect 8372 16044 9996 16100
rect 10052 16044 13804 16100
rect 13860 16044 13870 16100
rect 14018 16044 14028 16100
rect 14084 16044 16380 16100
rect 16436 16044 18508 16100
rect 18564 16044 18574 16100
rect 12114 15932 12124 15988
rect 12180 15932 14476 15988
rect 14532 15932 14542 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 20066 15260 20076 15316
rect 20132 15260 23324 15316
rect 23380 15260 25340 15316
rect 25396 15260 27132 15316
rect 27188 15260 28588 15316
rect 28644 15260 30044 15316
rect 30100 15260 30110 15316
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 14690 14700 14700 14756
rect 14756 14700 15708 14756
rect 15764 14700 15774 14756
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 25554 4060 25564 4116
rect 25620 4060 26796 4116
rect 26852 4060 26862 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 23538 3612 23548 3668
rect 23604 3612 24780 3668
rect 24836 3612 24846 3668
rect 16818 3388 16828 3444
rect 16884 3388 18060 3444
rect 18116 3388 18126 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 18060 21980 18116 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 18060 21196 18116 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 18060 22036 18116 22046
rect 18060 21252 18116 21980
rect 18060 21186 18116 21196
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18592 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22736 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _098_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21840 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _100_
timestamp 1698175906
transform -1 0 20944 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23408 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_
timestamp 1698175906
transform 1 0 18928 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1698175906
transform 1 0 17248 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform 1 0 22736 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26880 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 25984 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform -1 0 20944 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform -1 0 18816 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _110_
timestamp 1698175906
transform 1 0 18928 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform -1 0 20272 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform -1 0 21840 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _113_
timestamp 1698175906
transform -1 0 18816 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 18256 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20608 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20160 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22288 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _120_
timestamp 1698175906
transform 1 0 22288 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _121_
timestamp 1698175906
transform 1 0 22960 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _122_
timestamp 1698175906
transform -1 0 18592 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 19040 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 17472 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _125_
timestamp 1698175906
transform -1 0 14224 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _126_
timestamp 1698175906
transform 1 0 14224 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform -1 0 22960 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _128_
timestamp 1698175906
transform 1 0 16576 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform -1 0 14896 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14560 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 17920 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _133_
timestamp 1698175906
transform -1 0 14336 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1698175906
transform -1 0 19712 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform 1 0 19712 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _136_
timestamp 1698175906
transform -1 0 22848 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _137_
timestamp 1698175906
transform 1 0 20608 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform 1 0 18592 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform -1 0 20944 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform 1 0 17584 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _141_
timestamp 1698175906
transform -1 0 16576 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _143_
timestamp 1698175906
transform 1 0 13664 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16240 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1698175906
transform -1 0 16016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23184 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform -1 0 25760 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698175906
transform -1 0 16800 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _151_
timestamp 1698175906
transform -1 0 15680 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _152_
timestamp 1698175906
transform -1 0 20384 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform -1 0 15456 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _154_
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _155_
timestamp 1698175906
transform -1 0 19600 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _156_
timestamp 1698175906
transform -1 0 16576 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15344 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _158_
timestamp 1698175906
transform -1 0 13888 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform -1 0 12880 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _160_
timestamp 1698175906
transform 1 0 19600 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform -1 0 21728 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _162_
timestamp 1698175906
transform -1 0 20496 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform 1 0 21056 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 18816
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1698175906
transform 1 0 23296 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _168_
timestamp 1698175906
transform -1 0 23520 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 22512 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _170_
timestamp 1698175906
transform -1 0 16352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _171_
timestamp 1698175906
transform 1 0 16128 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform -1 0 15568 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 13104 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _174_
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _175_
timestamp 1698175906
transform 1 0 23408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform 1 0 28224 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _177_
timestamp 1698175906
transform -1 0 28224 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform 1 0 24304 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _179_
timestamp 1698175906
transform 1 0 25648 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _180_
timestamp 1698175906
transform -1 0 23408 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _182_
timestamp 1698175906
transform -1 0 26768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 25312 0 1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _185_
timestamp 1698175906
transform 1 0 26768 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _186_
timestamp 1698175906
transform -1 0 25760 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _187_
timestamp 1698175906
transform -1 0 24864 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _188_
timestamp 1698175906
transform -1 0 26320 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _189_
timestamp 1698175906
transform -1 0 25984 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform 1 0 16464 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform -1 0 13104 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform -1 0 13104 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform 1 0 19040 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 17696 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 19824 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform -1 0 14000 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 13776 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform -1 0 16128 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform -1 0 13104 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform -1 0 16800 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform -1 0 13104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 18704 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _205_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22736 0 1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 21280 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 13664 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform -1 0 13440 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 26768 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 26432 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 26768 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 23856 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 24864 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _218_
timestamp 1698175906
transform -1 0 26880 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _219_
timestamp 1698175906
transform 1 0 27104 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__CLK
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 23184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform -1 0 17696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 23296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 16128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 14112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 18480 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 27104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 24752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 14448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 30240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 29904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 30240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 28336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 17472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 23184 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698175906
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_243
timestamp 1698175906
transform 1 0 28560 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698175906
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698175906
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_131 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_139
timestamp 1698175906
transform 1 0 16912 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_143
timestamp 1698175906
transform 1 0 17360 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_107
timestamp 1698175906
transform 1 0 13328 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_162
timestamp 1698175906
transform 1 0 19488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_164
timestamp 1698175906
transform 1 0 19712 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_194
timestamp 1698175906
transform 1 0 23072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_198
timestamp 1698175906
transform 1 0 23520 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_241
timestamp 1698175906
transform 1 0 28336 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_245
timestamp 1698175906
transform 1 0 28784 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_69
timestamp 1698175906
transform 1 0 9072 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_73
timestamp 1698175906
transform 1 0 9520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_75
timestamp 1698175906
transform 1 0 9744 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_121
timestamp 1698175906
transform 1 0 14896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_129
timestamp 1698175906
transform 1 0 15792 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_143
timestamp 1698175906
transform 1 0 17360 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_228
timestamp 1698175906
transform 1 0 26880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_232
timestamp 1698175906
transform 1 0 27328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_240
timestamp 1698175906
transform 1 0 28224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_76
timestamp 1698175906
transform 1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_78
timestamp 1698175906
transform 1 0 10080 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698175906
transform 1 0 13440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698175906
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_169
timestamp 1698175906
transform 1 0 20272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_171
timestamp 1698175906
transform 1 0 20496 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_180
timestamp 1698175906
transform 1 0 21504 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_202
timestamp 1698175906
transform 1 0 23968 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_224
timestamp 1698175906
transform 1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_226
timestamp 1698175906
transform 1 0 26656 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_256
timestamp 1698175906
transform 1 0 30016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_260
timestamp 1698175906
transform 1 0 30464 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_85
timestamp 1698175906
transform 1 0 10864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_93
timestamp 1698175906
transform 1 0 11760 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_97
timestamp 1698175906
transform 1 0 12208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_99
timestamp 1698175906
transform 1 0 12432 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_119
timestamp 1698175906
transform 1 0 14672 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_135
timestamp 1698175906
transform 1 0 16464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_139
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_158
timestamp 1698175906
transform 1 0 19040 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_166
timestamp 1698175906
transform 1 0 19936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_170
timestamp 1698175906
transform 1 0 20384 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_211
timestamp 1698175906
transform 1 0 24976 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_219
timestamp 1698175906
transform 1 0 25872 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_228
timestamp 1698175906
transform 1 0 26880 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_120
timestamp 1698175906
transform 1 0 14784 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_128
timestamp 1698175906
transform 1 0 15680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_148
timestamp 1698175906
transform 1 0 17920 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_175
timestamp 1698175906
transform 1 0 20944 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_181
timestamp 1698175906
transform 1 0 21616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_228
timestamp 1698175906
transform 1 0 26880 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_232
timestamp 1698175906
transform 1 0 27328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_246
timestamp 1698175906
transform 1 0 28896 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_128
timestamp 1698175906
transform 1 0 15680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_134
timestamp 1698175906
transform 1 0 16352 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_144
timestamp 1698175906
transform 1 0 17472 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_192
timestamp 1698175906
transform 1 0 22848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_194
timestamp 1698175906
transform 1 0 23072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_215
timestamp 1698175906
transform 1 0 25424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_224
timestamp 1698175906
transform 1 0 26432 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_226
timestamp 1698175906
transform 1 0 26656 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_235
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 4480 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 8064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_96
timestamp 1698175906
transform 1 0 12096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698175906
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_170
timestamp 1698175906
transform 1 0 20384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_172
timestamp 1698175906
transform 1 0 20608 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_183
timestamp 1698175906
transform 1 0 21840 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_220
timestamp 1698175906
transform 1 0 25984 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_253
timestamp 1698175906
transform 1 0 29680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_257
timestamp 1698175906
transform 1 0 30128 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698175906
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 9744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_121
timestamp 1698175906
transform 1 0 14896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_194
timestamp 1698175906
transform 1 0 23072 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_253
timestamp 1698175906
transform 1 0 29680 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_285
timestamp 1698175906
transform 1 0 33264 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_301
timestamp 1698175906
transform 1 0 35056 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698175906
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698175906
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_112
timestamp 1698175906
transform 1 0 13888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_116
timestamp 1698175906
transform 1 0 14336 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_120
timestamp 1698175906
transform 1 0 14784 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_126
timestamp 1698175906
transform 1 0 15456 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_134
timestamp 1698175906
transform 1 0 16352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_218
timestamp 1698175906
transform 1 0 25760 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_256
timestamp 1698175906
transform 1 0 30016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_260
timestamp 1698175906
transform 1 0 30464 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_123
timestamp 1698175906
transform 1 0 15120 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_127
timestamp 1698175906
transform 1 0 15568 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_223
timestamp 1698175906
transform 1 0 26320 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_239
timestamp 1698175906
transform 1 0 28112 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_108
timestamp 1698175906
transform 1 0 13440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_118
timestamp 1698175906
transform 1 0 14560 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_122
timestamp 1698175906
transform 1 0 15008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_124
timestamp 1698175906
transform 1 0 15232 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_135
timestamp 1698175906
transform 1 0 16464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_148
timestamp 1698175906
transform 1 0 17920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_156
timestamp 1698175906
transform 1 0 18816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698175906
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_220
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_252
timestamp 1698175906
transform 1 0 29568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_268
timestamp 1698175906
transform 1 0 31360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_85
timestamp 1698175906
transform 1 0 10864 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698175906
transform 1 0 11760 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_97
timestamp 1698175906
transform 1 0 12208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_138
timestamp 1698175906
transform 1 0 16800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_142
timestamp 1698175906
transform 1 0 17248 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_150
timestamp 1698175906
transform 1 0 18144 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_154
timestamp 1698175906
transform 1 0 18592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_156
timestamp 1698175906
transform 1 0 18816 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_164
timestamp 1698175906
transform 1 0 19712 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_168
timestamp 1698175906
transform 1 0 20160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_193
timestamp 1698175906
transform 1 0 22960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_197
timestamp 1698175906
transform 1 0 23408 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_239
timestamp 1698175906
transform 1 0 28112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_118
timestamp 1698175906
transform 1 0 14560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_122
timestamp 1698175906
transform 1 0 15008 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698175906
transform 1 0 16352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_158
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_162
timestamp 1698175906
transform 1 0 19488 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_171
timestamp 1698175906
transform 1 0 20496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_175
timestamp 1698175906
transform 1 0 20944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_183
timestamp 1698175906
transform 1 0 21840 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_199
timestamp 1698175906
transform 1 0 23632 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698175906
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_218
timestamp 1698175906
transform 1 0 25760 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_250
timestamp 1698175906
transform 1 0 29344 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698175906
transform 1 0 31136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_69
timestamp 1698175906
transform 1 0 9072 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_73
timestamp 1698175906
transform 1 0 9520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_75
timestamp 1698175906
transform 1 0 9744 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_116
timestamp 1698175906
transform 1 0 14336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_120
timestamp 1698175906
transform 1 0 14784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_127
timestamp 1698175906
transform 1 0 15568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_131
timestamp 1698175906
transform 1 0 16016 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_140
timestamp 1698175906
transform 1 0 17024 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_148
timestamp 1698175906
transform 1 0 17920 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_152
timestamp 1698175906
transform 1 0 18368 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_155
timestamp 1698175906
transform 1 0 18704 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1698175906
transform 1 0 20160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_182
timestamp 1698175906
transform 1 0 21728 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_198
timestamp 1698175906
transform 1 0 23520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_200
timestamp 1698175906
transform 1 0 23744 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_236
timestamp 1698175906
transform 1 0 27776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698175906
transform 1 0 28224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_107
timestamp 1698175906
transform 1 0 13328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_109
timestamp 1698175906
transform 1 0 13552 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_198
timestamp 1698175906
transform 1 0 23520 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_131
timestamp 1698175906
transform 1 0 16016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_207
timestamp 1698175906
transform 1 0 24528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_211
timestamp 1698175906
transform 1 0 24976 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_333
timestamp 1698175906
transform 1 0 38640 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_341
timestamp 1698175906
transform 1 0 39536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698175906
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_341
timestamp 1698175906
transform 1 0 39536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698175906
transform 1 0 19040 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_189
timestamp 1698175906
transform 1 0 22512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698175906
transform 1 0 24304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 20272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita3_23 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39984 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita3_24
timestamp 1698175906
transform 1 0 39984 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita3_25
timestamp 1698175906
transform -1 0 20272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita3_26
timestamp 1698175906
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 16912 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 25648 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 27328 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 4480 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 4480 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 16912 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 19600 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 36288 42000 36400 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 21504 41200 21616 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 18816 41200 18928 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 26488 20776 26488 20776 0 _000_
rlabel metal2 27720 20804 27720 20804 0 _001_
rlabel metal2 24360 24696 24360 24696 0 _002_
rlabel metal2 25704 23576 25704 23576 0 _003_
rlabel metal2 26040 16072 26040 16072 0 _004_
rlabel metal2 17752 26936 17752 26936 0 _005_
rlabel metal3 13328 15960 13328 15960 0 _006_
rlabel metal3 13104 25368 13104 25368 0 _007_
rlabel metal2 19824 20104 19824 20104 0 _008_
rlabel metal2 18648 14868 18648 14868 0 _009_
rlabel metal2 20832 15400 20832 15400 0 _010_
rlabel metal2 14728 17584 14728 17584 0 _011_
rlabel metal2 12824 24304 12824 24304 0 _012_
rlabel metal3 15232 14728 15232 14728 0 _013_
rlabel metal2 15176 19656 15176 19656 0 _014_
rlabel metal2 13496 20552 13496 20552 0 _015_
rlabel metal2 15848 23576 15848 23576 0 _016_
rlabel metal2 12376 20440 12376 20440 0 _017_
rlabel metal2 19712 26824 19712 26824 0 _018_
rlabel metal2 23688 16464 23688 16464 0 _019_
rlabel metal2 22120 26936 22120 26936 0 _020_
rlabel metal2 15064 25816 15064 25816 0 _021_
rlabel metal2 12488 17192 12488 17192 0 _022_
rlabel metal2 27720 17584 27720 17584 0 _023_
rlabel metal2 15848 14840 15848 14840 0 _024_
rlabel metal2 25592 21952 25592 21952 0 _025_
rlabel metal2 15960 22736 15960 22736 0 _026_
rlabel metal2 15568 19208 15568 19208 0 _027_
rlabel metal2 13832 18648 13832 18648 0 _028_
rlabel metal2 13552 20776 13552 20776 0 _029_
rlabel metal2 16520 21056 16520 21056 0 _030_
rlabel metal2 16296 22792 16296 22792 0 _031_
rlabel metal2 13104 21336 13104 21336 0 _032_
rlabel metal3 21056 26936 21056 26936 0 _033_
rlabel metal2 20832 27048 20832 27048 0 _034_
rlabel metal3 21952 18424 21952 18424 0 _035_
rlabel metal2 23464 17528 23464 17528 0 _036_
rlabel metal2 23128 24864 23128 24864 0 _037_
rlabel metal2 25368 22680 25368 22680 0 _038_
rlabel metal2 22344 26432 22344 26432 0 _039_
rlabel metal2 16072 24976 16072 24976 0 _040_
rlabel metal2 15904 25480 15904 25480 0 _041_
rlabel metal3 12992 17640 12992 17640 0 _042_
rlabel metal2 27720 19096 27720 19096 0 _043_
rlabel metal2 28280 18424 28280 18424 0 _044_
rlabel metal2 24808 20832 24808 20832 0 _045_
rlabel metal2 26376 19656 26376 19656 0 _046_
rlabel metal2 22904 20496 22904 20496 0 _047_
rlabel metal2 27328 19432 27328 19432 0 _048_
rlabel metal3 28224 20552 28224 20552 0 _049_
rlabel metal2 27048 20720 27048 20720 0 _050_
rlabel metal2 24696 24192 24696 24192 0 _051_
rlabel metal2 25816 22792 25816 22792 0 _052_
rlabel metal2 18648 18816 18648 18816 0 _053_
rlabel metal2 24080 17640 24080 17640 0 _054_
rlabel metal3 18200 18424 18200 18424 0 _055_
rlabel metal2 25032 19992 25032 19992 0 _056_
rlabel metal2 19544 21168 19544 21168 0 _057_
rlabel metal3 18592 16856 18592 16856 0 _058_
rlabel metal2 24808 17248 24808 17248 0 _059_
rlabel metal2 19208 18984 19208 18984 0 _060_
rlabel metal2 28392 17696 28392 17696 0 _061_
rlabel metal2 14840 18256 14840 18256 0 _062_
rlabel metal3 23576 18536 23576 18536 0 _063_
rlabel metal2 25816 17024 25816 17024 0 _064_
rlabel metal2 18872 21504 18872 21504 0 _065_
rlabel metal3 17024 23240 17024 23240 0 _066_
rlabel metal3 21616 18312 21616 18312 0 _067_
rlabel metal2 19768 19320 19768 19320 0 _068_
rlabel metal2 20664 23632 20664 23632 0 _069_
rlabel metal2 18032 22344 18032 22344 0 _070_
rlabel metal2 18984 20188 18984 20188 0 _071_
rlabel metal2 19712 25256 19712 25256 0 _072_
rlabel metal2 19432 25928 19432 25928 0 _073_
rlabel metal2 17864 21392 17864 21392 0 _074_
rlabel metal3 19824 22232 19824 22232 0 _075_
rlabel metal2 23128 22008 23128 22008 0 _076_
rlabel metal2 24024 23240 24024 23240 0 _077_
rlabel metal2 15064 17640 15064 17640 0 _078_
rlabel metal2 13944 17136 13944 17136 0 _079_
rlabel metal2 13720 20860 13720 20860 0 _080_
rlabel metal2 13944 15736 13944 15736 0 _081_
rlabel metal3 19880 19096 19880 19096 0 _082_
rlabel metal2 13832 25592 13832 25592 0 _083_
rlabel metal2 13832 23800 13832 23800 0 _084_
rlabel metal2 14112 24920 14112 24920 0 _085_
rlabel metal2 13720 25368 13720 25368 0 _086_
rlabel metal2 20440 16856 20440 16856 0 _087_
rlabel metal2 21840 19320 21840 19320 0 _088_
rlabel metal3 19936 21784 19936 21784 0 _089_
rlabel metal2 20440 22904 20440 22904 0 _090_
rlabel metal2 16408 18704 16408 18704 0 _091_
rlabel metal2 14392 22512 14392 22512 0 _092_
rlabel metal3 13440 23352 13440 23352 0 _093_
rlabel metal2 17192 16184 17192 16184 0 _094_
rlabel metal3 2478 26936 2478 26936 0 clk
rlabel metal2 23352 21112 23352 21112 0 clknet_0_clk
rlabel metal2 13944 25424 13944 25424 0 clknet_1_0__leaf_clk
rlabel metal3 23184 27048 23184 27048 0 clknet_1_1__leaf_clk
rlabel metal2 21560 19992 21560 19992 0 dut3.count\[0\]
rlabel metal2 20888 14616 20888 14616 0 dut3.count\[1\]
rlabel metal2 22568 16296 22568 16296 0 dut3.count\[2\]
rlabel metal3 18088 17528 18088 17528 0 dut3.count\[3\]
rlabel metal2 29512 19488 29512 19488 0 net1
rlabel metal2 37912 25760 37912 25760 0 net10
rlabel metal3 6356 20776 6356 20776 0 net11
rlabel metal2 10360 17192 10360 17192 0 net12
rlabel metal2 29848 17584 29848 17584 0 net13
rlabel metal2 13720 23968 13720 23968 0 net14
rlabel metal3 6356 21560 6356 21560 0 net15
rlabel metal2 13048 19936 13048 19936 0 net16
rlabel metal2 17080 5964 17080 5964 0 net17
rlabel metal3 6356 24696 6356 24696 0 net18
rlabel metal3 6356 25480 6356 25480 0 net19
rlabel metal2 27384 25536 27384 25536 0 net2
rlabel metal2 4312 16576 4312 16576 0 net20
rlabel metal2 28168 16408 28168 16408 0 net21
rlabel metal2 19656 37240 19656 37240 0 net22
rlabel metal2 40264 26544 40264 26544 0 net23
rlabel metal3 40754 36344 40754 36344 0 net24
rlabel metal2 19992 38248 19992 38248 0 net25
rlabel metal3 1246 36344 1246 36344 0 net26
rlabel metal2 24360 29540 24360 29540 0 net3
rlabel metal2 16744 26208 16744 26208 0 net4
rlabel metal2 27944 23576 27944 23576 0 net5
rlabel metal2 21784 26096 21784 26096 0 net6
rlabel metal2 25816 6356 25816 6356 0 net7
rlabel metal2 27160 5964 27160 5964 0 net8
rlabel metal2 29512 20664 29512 20664 0 net9
rlabel metal2 39928 21168 39928 21168 0 segm[0]
rlabel metal2 40040 25256 40040 25256 0 segm[10]
rlabel metal2 24248 39746 24248 39746 0 segm[11]
rlabel metal2 16856 39746 16856 39746 0 segm[12]
rlabel metal3 40642 22904 40642 22904 0 segm[13]
rlabel metal2 21560 39746 21560 39746 0 segm[3]
rlabel metal2 25592 2422 25592 2422 0 segm[6]
rlabel metal2 23576 2198 23576 2198 0 segm[7]
rlabel metal2 40040 20552 40040 20552 0 segm[8]
rlabel metal2 39928 25872 39928 25872 0 segm[9]
rlabel metal3 1414 20216 1414 20216 0 sel[0]
rlabel metal3 1358 16856 1358 16856 0 sel[10]
rlabel metal3 40642 18200 40642 18200 0 sel[11]
rlabel metal3 1358 23576 1358 23576 0 sel[1]
rlabel metal3 1358 20888 1358 20888 0 sel[2]
rlabel metal3 1358 19544 1358 19544 0 sel[3]
rlabel metal2 16856 2086 16856 2086 0 sel[4]
rlabel metal3 1358 24248 1358 24248 0 sel[5]
rlabel metal3 1358 24920 1358 24920 0 sel[6]
rlabel metal3 1358 16184 1358 16184 0 sel[7]
rlabel metal2 40040 17304 40040 17304 0 sel[8]
rlabel metal2 19544 39354 19544 39354 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
