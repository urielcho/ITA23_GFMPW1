magic
tech gf180mcuD
magscale 1 10
timestamp 1699641377
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 22430 38274 22482 38286
rect 19506 38222 19518 38274
rect 19570 38222 19582 38274
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 14802 38110 14814 38162
rect 14866 38110 14878 38162
rect 15922 37998 15934 38050
rect 15986 37998 15998 38050
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 21410 37998 21422 38050
rect 21474 37998 21486 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 1710 37378 1762 37390
rect 1710 37314 1762 37326
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 20850 37214 20862 37266
rect 20914 37214 20926 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 16718 36706 16770 36718
rect 16718 36642 16770 36654
rect 15698 36430 15710 36482
rect 15762 36430 15774 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 13458 28702 13470 28754
rect 13522 28702 13534 28754
rect 16830 28642 16882 28654
rect 16258 28590 16270 28642
rect 16322 28590 16334 28642
rect 16830 28578 16882 28590
rect 18510 28530 18562 28542
rect 15586 28478 15598 28530
rect 15650 28478 15662 28530
rect 18510 28466 18562 28478
rect 18622 28530 18674 28542
rect 18622 28466 18674 28478
rect 18846 28418 18898 28430
rect 18846 28354 18898 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 14926 28082 14978 28094
rect 15486 28082 15538 28094
rect 15250 28030 15262 28082
rect 15314 28030 15326 28082
rect 14926 28018 14978 28030
rect 15486 28018 15538 28030
rect 15710 27970 15762 27982
rect 15710 27906 15762 27918
rect 15822 27858 15874 27870
rect 14130 27806 14142 27858
rect 14194 27806 14206 27858
rect 20290 27806 20302 27858
rect 20354 27806 20366 27858
rect 15822 27794 15874 27806
rect 14590 27746 14642 27758
rect 20750 27746 20802 27758
rect 11218 27694 11230 27746
rect 11282 27694 11294 27746
rect 13346 27694 13358 27746
rect 13410 27694 13422 27746
rect 17378 27694 17390 27746
rect 17442 27694 17454 27746
rect 19506 27694 19518 27746
rect 19570 27694 19582 27746
rect 14590 27682 14642 27694
rect 20750 27682 20802 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 15598 27298 15650 27310
rect 15598 27234 15650 27246
rect 1934 27186 1986 27198
rect 1934 27122 1986 27134
rect 13918 27074 13970 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 13918 27010 13970 27022
rect 15150 27074 15202 27086
rect 15150 27010 15202 27022
rect 19070 27074 19122 27086
rect 19070 27010 19122 27022
rect 19406 27074 19458 27086
rect 19406 27010 19458 27022
rect 13806 26962 13858 26974
rect 13806 26898 13858 26910
rect 14254 26962 14306 26974
rect 14254 26898 14306 26910
rect 14590 26962 14642 26974
rect 14590 26898 14642 26910
rect 14814 26962 14866 26974
rect 14814 26898 14866 26910
rect 15038 26962 15090 26974
rect 15038 26898 15090 26910
rect 15598 26962 15650 26974
rect 15598 26898 15650 26910
rect 15710 26962 15762 26974
rect 15710 26898 15762 26910
rect 21870 26962 21922 26974
rect 21870 26898 21922 26910
rect 22094 26962 22146 26974
rect 22094 26898 22146 26910
rect 22206 26962 22258 26974
rect 22206 26898 22258 26910
rect 13582 26850 13634 26862
rect 13582 26786 13634 26798
rect 14478 26850 14530 26862
rect 14478 26786 14530 26798
rect 19182 26850 19234 26862
rect 19182 26786 19234 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 17938 26462 17950 26514
rect 18002 26462 18014 26514
rect 13122 26350 13134 26402
rect 13186 26350 13198 26402
rect 25554 26350 25566 26402
rect 25618 26350 25630 26402
rect 12450 26238 12462 26290
rect 12514 26238 12526 26290
rect 18162 26238 18174 26290
rect 18226 26238 18238 26290
rect 20402 26238 20414 26290
rect 20466 26238 20478 26290
rect 25330 26238 25342 26290
rect 25394 26238 25406 26290
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 15710 26178 15762 26190
rect 15250 26126 15262 26178
rect 15314 26126 15326 26178
rect 15710 26114 15762 26126
rect 19518 26178 19570 26190
rect 19518 26114 19570 26126
rect 19966 26178 20018 26190
rect 21074 26126 21086 26178
rect 21138 26126 21150 26178
rect 23202 26126 23214 26178
rect 23266 26126 23278 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 19966 26114 20018 26126
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 13918 25730 13970 25742
rect 13918 25666 13970 25678
rect 21310 25730 21362 25742
rect 21310 25666 21362 25678
rect 21422 25730 21474 25742
rect 21422 25666 21474 25678
rect 40014 25618 40066 25630
rect 20626 25566 20638 25618
rect 20690 25566 20702 25618
rect 40014 25554 40066 25566
rect 13694 25506 13746 25518
rect 21870 25506 21922 25518
rect 17714 25454 17726 25506
rect 17778 25454 17790 25506
rect 13694 25442 13746 25454
rect 21870 25442 21922 25454
rect 22094 25506 22146 25518
rect 22754 25454 22766 25506
rect 22818 25454 22830 25506
rect 37874 25454 37886 25506
rect 37938 25454 37950 25506
rect 22094 25442 22146 25454
rect 14254 25394 14306 25406
rect 14254 25330 14306 25342
rect 15374 25394 15426 25406
rect 21534 25394 21586 25406
rect 18498 25342 18510 25394
rect 18562 25342 18574 25394
rect 23538 25342 23550 25394
rect 23602 25342 23614 25394
rect 15374 25330 15426 25342
rect 21534 25330 21586 25342
rect 14030 25282 14082 25294
rect 14030 25218 14082 25230
rect 14926 25282 14978 25294
rect 14926 25218 14978 25230
rect 15038 25282 15090 25294
rect 15038 25218 15090 25230
rect 15150 25282 15202 25294
rect 26238 25282 26290 25294
rect 25778 25230 25790 25282
rect 25842 25230 25854 25282
rect 26562 25230 26574 25282
rect 26626 25230 26638 25282
rect 15150 25218 15202 25230
rect 26238 25218 26290 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 13470 24946 13522 24958
rect 13470 24882 13522 24894
rect 13694 24946 13746 24958
rect 13694 24882 13746 24894
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 23774 24946 23826 24958
rect 23774 24882 23826 24894
rect 14690 24782 14702 24834
rect 14754 24782 14766 24834
rect 18274 24782 18286 24834
rect 18338 24782 18350 24834
rect 13358 24722 13410 24734
rect 24670 24722 24722 24734
rect 14018 24670 14030 24722
rect 14082 24670 14094 24722
rect 23314 24670 23326 24722
rect 23378 24670 23390 24722
rect 23986 24670 23998 24722
rect 24050 24670 24062 24722
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 13358 24658 13410 24670
rect 24670 24658 24722 24670
rect 16818 24558 16830 24610
rect 16882 24558 16894 24610
rect 26002 24558 26014 24610
rect 26066 24558 26078 24610
rect 28130 24558 28142 24610
rect 28194 24558 28206 24610
rect 23662 24498 23714 24510
rect 23662 24434 23714 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 18174 24162 18226 24174
rect 18174 24098 18226 24110
rect 13694 24050 13746 24062
rect 22430 24050 22482 24062
rect 19394 23998 19406 24050
rect 19458 23998 19470 24050
rect 13694 23986 13746 23998
rect 22430 23986 22482 23998
rect 25230 24050 25282 24062
rect 25230 23986 25282 23998
rect 40014 24050 40066 24062
rect 40014 23986 40066 23998
rect 13806 23938 13858 23950
rect 19630 23938 19682 23950
rect 14354 23886 14366 23938
rect 14418 23886 14430 23938
rect 17266 23886 17278 23938
rect 17330 23886 17342 23938
rect 13806 23874 13858 23886
rect 19630 23874 19682 23886
rect 20078 23938 20130 23950
rect 20078 23874 20130 23886
rect 20190 23938 20242 23950
rect 20190 23874 20242 23886
rect 22766 23938 22818 23950
rect 22766 23874 22818 23886
rect 23774 23938 23826 23950
rect 23774 23874 23826 23886
rect 23886 23938 23938 23950
rect 23886 23874 23938 23886
rect 25118 23938 25170 23950
rect 25118 23874 25170 23886
rect 25790 23938 25842 23950
rect 25790 23874 25842 23886
rect 26126 23938 26178 23950
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 26126 23874 26178 23886
rect 17838 23826 17890 23838
rect 17838 23762 17890 23774
rect 19406 23826 19458 23838
rect 23438 23826 23490 23838
rect 23090 23774 23102 23826
rect 23154 23774 23166 23826
rect 19406 23762 19458 23774
rect 23438 23762 23490 23774
rect 26350 23826 26402 23838
rect 26350 23762 26402 23774
rect 26462 23826 26514 23838
rect 26462 23762 26514 23774
rect 18062 23714 18114 23726
rect 17490 23662 17502 23714
rect 17554 23662 17566 23714
rect 18062 23650 18114 23662
rect 19966 23714 20018 23726
rect 19966 23650 20018 23662
rect 20414 23714 20466 23726
rect 20414 23650 20466 23662
rect 23662 23714 23714 23726
rect 23662 23650 23714 23662
rect 25342 23714 25394 23726
rect 25342 23650 25394 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 15374 23378 15426 23390
rect 15374 23314 15426 23326
rect 22766 23378 22818 23390
rect 22766 23314 22818 23326
rect 14142 23266 14194 23278
rect 14142 23202 14194 23214
rect 14366 23266 14418 23278
rect 14366 23202 14418 23214
rect 15150 23266 15202 23278
rect 15150 23202 15202 23214
rect 15598 23266 15650 23278
rect 15598 23202 15650 23214
rect 15710 23154 15762 23166
rect 10994 23102 11006 23154
rect 11058 23102 11070 23154
rect 14914 23102 14926 23154
rect 14978 23102 14990 23154
rect 19394 23102 19406 23154
rect 19458 23102 19470 23154
rect 15710 23090 15762 23102
rect 14254 23042 14306 23054
rect 11666 22990 11678 23042
rect 11730 22990 11742 23042
rect 13794 22990 13806 23042
rect 13858 22990 13870 23042
rect 14254 22978 14306 22990
rect 17502 23042 17554 23054
rect 20178 22990 20190 23042
rect 20242 22990 20254 23042
rect 22306 22990 22318 23042
rect 22370 22990 22382 23042
rect 17502 22978 17554 22990
rect 17614 22930 17666 22942
rect 17614 22866 17666 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 14478 22594 14530 22606
rect 14478 22530 14530 22542
rect 15038 22594 15090 22606
rect 15038 22530 15090 22542
rect 15822 22594 15874 22606
rect 15822 22530 15874 22542
rect 24894 22482 24946 22494
rect 24894 22418 24946 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 14926 22370 14978 22382
rect 22766 22370 22818 22382
rect 16146 22318 16158 22370
rect 16210 22318 16222 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 14926 22306 14978 22318
rect 22766 22306 22818 22318
rect 14590 22258 14642 22270
rect 14590 22194 14642 22206
rect 15934 22258 15986 22270
rect 15934 22194 15986 22206
rect 17390 22258 17442 22270
rect 17390 22194 17442 22206
rect 17614 22258 17666 22270
rect 17614 22194 17666 22206
rect 19630 22258 19682 22270
rect 19630 22194 19682 22206
rect 19742 22258 19794 22270
rect 19742 22194 19794 22206
rect 19966 22258 20018 22270
rect 19966 22194 20018 22206
rect 21422 22258 21474 22270
rect 21422 22194 21474 22206
rect 21534 22258 21586 22270
rect 21534 22194 21586 22206
rect 22430 22258 22482 22270
rect 22430 22194 22482 22206
rect 22542 22258 22594 22270
rect 22542 22194 22594 22206
rect 14030 22146 14082 22158
rect 14030 22082 14082 22094
rect 14478 22146 14530 22158
rect 14478 22082 14530 22094
rect 17502 22146 17554 22158
rect 17502 22082 17554 22094
rect 18174 22146 18226 22158
rect 18958 22146 19010 22158
rect 18498 22094 18510 22146
rect 18562 22094 18574 22146
rect 18174 22082 18226 22094
rect 18958 22082 19010 22094
rect 20190 22146 20242 22158
rect 21198 22146 21250 22158
rect 20514 22094 20526 22146
rect 20578 22094 20590 22146
rect 20190 22082 20242 22094
rect 21198 22082 21250 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14590 21810 14642 21822
rect 24322 21758 24334 21810
rect 24386 21758 24398 21810
rect 14590 21746 14642 21758
rect 14914 21646 14926 21698
rect 14978 21646 14990 21698
rect 28802 21646 28814 21698
rect 28866 21646 28878 21698
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 18610 21534 18622 21586
rect 18674 21534 18686 21586
rect 24098 21534 24110 21586
rect 24162 21534 24174 21586
rect 25218 21534 25230 21586
rect 25282 21534 25294 21586
rect 28578 21534 28590 21586
rect 28642 21534 28654 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 13134 21474 13186 21486
rect 13134 21410 13186 21422
rect 17502 21474 17554 21486
rect 17502 21410 17554 21422
rect 17726 21474 17778 21486
rect 40014 21474 40066 21486
rect 23426 21422 23438 21474
rect 23490 21422 23502 21474
rect 26002 21422 26014 21474
rect 26066 21422 26078 21474
rect 28130 21422 28142 21474
rect 28194 21422 28206 21474
rect 17726 21410 17778 21422
rect 40014 21410 40066 21422
rect 1934 21362 1986 21374
rect 1934 21298 1986 21310
rect 18062 21362 18114 21374
rect 18062 21298 18114 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 13918 21026 13970 21038
rect 13918 20962 13970 20974
rect 15038 21026 15090 21038
rect 24222 21026 24274 21038
rect 17938 20974 17950 21026
rect 18002 20974 18014 21026
rect 15038 20962 15090 20974
rect 24222 20962 24274 20974
rect 19966 20914 20018 20926
rect 9986 20862 9998 20914
rect 10050 20862 10062 20914
rect 17154 20862 17166 20914
rect 17218 20862 17230 20914
rect 19966 20850 20018 20862
rect 23214 20914 23266 20926
rect 23214 20850 23266 20862
rect 24446 20914 24498 20926
rect 24446 20850 24498 20862
rect 24558 20914 24610 20926
rect 24558 20850 24610 20862
rect 27022 20914 27074 20926
rect 27022 20850 27074 20862
rect 40014 20914 40066 20926
rect 40014 20850 40066 20862
rect 14478 20802 14530 20814
rect 12898 20750 12910 20802
rect 12962 20750 12974 20802
rect 13570 20750 13582 20802
rect 13634 20750 13646 20802
rect 14478 20738 14530 20750
rect 14926 20802 14978 20814
rect 14926 20738 14978 20750
rect 15262 20802 15314 20814
rect 15262 20738 15314 20750
rect 16158 20802 16210 20814
rect 20078 20802 20130 20814
rect 17378 20750 17390 20802
rect 17442 20750 17454 20802
rect 17714 20750 17726 20802
rect 17778 20750 17790 20802
rect 19618 20750 19630 20802
rect 19682 20750 19694 20802
rect 16158 20738 16210 20750
rect 20078 20738 20130 20750
rect 21310 20802 21362 20814
rect 22194 20750 22206 20802
rect 22258 20750 22270 20802
rect 23762 20750 23774 20802
rect 23826 20750 23838 20802
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 21310 20738 21362 20750
rect 15374 20690 15426 20702
rect 12114 20638 12126 20690
rect 12178 20638 12190 20690
rect 15374 20626 15426 20638
rect 15486 20690 15538 20702
rect 19854 20690 19906 20702
rect 15810 20638 15822 20690
rect 15874 20638 15886 20690
rect 15486 20626 15538 20638
rect 19854 20626 19906 20638
rect 20302 20690 20354 20702
rect 20302 20626 20354 20638
rect 23102 20690 23154 20702
rect 24670 20690 24722 20702
rect 23986 20638 23998 20690
rect 24050 20638 24062 20690
rect 23102 20626 23154 20638
rect 24670 20626 24722 20638
rect 26014 20690 26066 20702
rect 26014 20626 26066 20638
rect 26910 20690 26962 20702
rect 26910 20626 26962 20638
rect 13806 20578 13858 20590
rect 13806 20514 13858 20526
rect 18846 20578 18898 20590
rect 23326 20578 23378 20590
rect 19170 20526 19182 20578
rect 19234 20526 19246 20578
rect 21634 20526 21646 20578
rect 21698 20526 21710 20578
rect 21970 20526 21982 20578
rect 22034 20526 22046 20578
rect 18846 20514 18898 20526
rect 23326 20514 23378 20526
rect 26126 20578 26178 20590
rect 26126 20514 26178 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 14478 20242 14530 20254
rect 14478 20178 14530 20190
rect 16382 20242 16434 20254
rect 16382 20178 16434 20190
rect 18622 20242 18674 20254
rect 18622 20178 18674 20190
rect 14702 20130 14754 20142
rect 12114 20078 12126 20130
rect 12178 20078 12190 20130
rect 14702 20066 14754 20078
rect 14814 20130 14866 20142
rect 14814 20066 14866 20078
rect 18062 20130 18114 20142
rect 18946 20078 18958 20130
rect 19010 20078 19022 20130
rect 20850 20078 20862 20130
rect 20914 20078 20926 20130
rect 26226 20078 26238 20130
rect 26290 20078 26302 20130
rect 18062 20066 18114 20078
rect 11442 19966 11454 20018
rect 11506 19966 11518 20018
rect 16258 19966 16270 20018
rect 16322 19966 16334 20018
rect 18274 19966 18286 20018
rect 18338 19966 18350 20018
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 20290 19966 20302 20018
rect 20354 19966 20366 20018
rect 25442 19966 25454 20018
rect 25506 19966 25518 20018
rect 15374 19906 15426 19918
rect 21422 19906 21474 19918
rect 14242 19854 14254 19906
rect 14306 19854 14318 19906
rect 16146 19854 16158 19906
rect 16210 19854 16222 19906
rect 20178 19854 20190 19906
rect 20242 19854 20254 19906
rect 15374 19842 15426 19854
rect 21422 19842 21474 19854
rect 24782 19906 24834 19918
rect 28354 19854 28366 19906
rect 28418 19854 28430 19906
rect 24782 19842 24834 19854
rect 17950 19794 18002 19806
rect 17950 19730 18002 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 17726 19458 17778 19470
rect 15810 19406 15822 19458
rect 15874 19406 15886 19458
rect 17726 19394 17778 19406
rect 15486 19346 15538 19358
rect 15486 19282 15538 19294
rect 16382 19346 16434 19358
rect 16382 19282 16434 19294
rect 17838 19346 17890 19358
rect 25454 19346 25506 19358
rect 19058 19294 19070 19346
rect 19122 19294 19134 19346
rect 22082 19294 22094 19346
rect 22146 19294 22158 19346
rect 24210 19294 24222 19346
rect 24274 19294 24286 19346
rect 17838 19282 17890 19294
rect 25454 19282 25506 19294
rect 14926 19234 14978 19246
rect 14926 19170 14978 19182
rect 16158 19234 16210 19246
rect 16158 19170 16210 19182
rect 17054 19234 17106 19246
rect 18958 19234 19010 19246
rect 18050 19182 18062 19234
rect 18114 19182 18126 19234
rect 19394 19182 19406 19234
rect 19458 19182 19470 19234
rect 21410 19182 21422 19234
rect 21474 19182 21486 19234
rect 25106 19182 25118 19234
rect 25170 19182 25182 19234
rect 25778 19182 25790 19234
rect 25842 19182 25854 19234
rect 17054 19170 17106 19182
rect 18958 19170 19010 19182
rect 20414 19122 20466 19134
rect 20414 19058 20466 19070
rect 25566 19122 25618 19134
rect 25566 19058 25618 19070
rect 25342 19010 25394 19022
rect 17378 18958 17390 19010
rect 17442 18958 17454 19010
rect 19954 18958 19966 19010
rect 20018 18958 20030 19010
rect 20738 18958 20750 19010
rect 20802 18958 20814 19010
rect 25342 18946 25394 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 18622 18674 18674 18686
rect 22318 18674 22370 18686
rect 25902 18674 25954 18686
rect 16818 18622 16830 18674
rect 16882 18622 16894 18674
rect 19170 18622 19182 18674
rect 19234 18622 19246 18674
rect 23538 18622 23550 18674
rect 23602 18622 23614 18674
rect 18622 18610 18674 18622
rect 22318 18610 22370 18622
rect 25902 18610 25954 18622
rect 18734 18562 18786 18574
rect 21870 18562 21922 18574
rect 17714 18510 17726 18562
rect 17778 18510 17790 18562
rect 19058 18510 19070 18562
rect 19122 18510 19134 18562
rect 20738 18510 20750 18562
rect 20802 18510 20814 18562
rect 18734 18498 18786 18510
rect 21870 18498 21922 18510
rect 22430 18562 22482 18574
rect 22430 18498 22482 18510
rect 16494 18450 16546 18462
rect 16494 18386 16546 18398
rect 18062 18450 18114 18462
rect 21982 18450 22034 18462
rect 25230 18450 25282 18462
rect 18386 18398 18398 18450
rect 18450 18398 18462 18450
rect 19618 18398 19630 18450
rect 19682 18398 19694 18450
rect 20066 18398 20078 18450
rect 20130 18398 20142 18450
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 23762 18398 23774 18450
rect 23826 18398 23838 18450
rect 18062 18386 18114 18398
rect 21982 18386 22034 18398
rect 25230 18386 25282 18398
rect 25678 18450 25730 18462
rect 25678 18386 25730 18398
rect 26126 18450 26178 18462
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 26126 18386 26178 18398
rect 25454 18338 25506 18350
rect 21298 18286 21310 18338
rect 21362 18286 21374 18338
rect 26002 18286 26014 18338
rect 26066 18286 26078 18338
rect 25454 18274 25506 18286
rect 21086 18226 21138 18238
rect 21086 18162 21138 18174
rect 21870 18226 21922 18238
rect 21870 18162 21922 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 17950 17890 18002 17902
rect 17950 17826 18002 17838
rect 18062 17890 18114 17902
rect 18062 17826 18114 17838
rect 18286 17890 18338 17902
rect 18286 17826 18338 17838
rect 18846 17890 18898 17902
rect 18846 17826 18898 17838
rect 19630 17890 19682 17902
rect 19630 17826 19682 17838
rect 20190 17890 20242 17902
rect 20190 17826 20242 17838
rect 20302 17890 20354 17902
rect 20302 17826 20354 17838
rect 21982 17890 22034 17902
rect 21982 17826 22034 17838
rect 22654 17890 22706 17902
rect 22654 17826 22706 17838
rect 1934 17778 1986 17790
rect 1934 17714 1986 17726
rect 15038 17778 15090 17790
rect 15038 17714 15090 17726
rect 21870 17778 21922 17790
rect 22978 17726 22990 17778
rect 23042 17726 23054 17778
rect 25890 17726 25902 17778
rect 25954 17726 25966 17778
rect 28018 17726 28030 17778
rect 28082 17726 28094 17778
rect 21870 17714 21922 17726
rect 14366 17666 14418 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 14366 17602 14418 17614
rect 14702 17666 14754 17678
rect 14702 17602 14754 17614
rect 15262 17666 15314 17678
rect 15262 17602 15314 17614
rect 15486 17666 15538 17678
rect 15486 17602 15538 17614
rect 17054 17666 17106 17678
rect 17054 17602 17106 17614
rect 18398 17666 18450 17678
rect 18398 17602 18450 17614
rect 19070 17666 19122 17678
rect 19070 17602 19122 17614
rect 19406 17666 19458 17678
rect 19406 17602 19458 17614
rect 20526 17666 20578 17678
rect 20526 17602 20578 17614
rect 21534 17666 21586 17678
rect 25106 17614 25118 17666
rect 25170 17614 25182 17666
rect 21534 17602 21586 17614
rect 14030 17554 14082 17566
rect 14030 17490 14082 17502
rect 14926 17554 14978 17566
rect 19182 17554 19234 17566
rect 17378 17502 17390 17554
rect 17442 17502 17454 17554
rect 14926 17490 14978 17502
rect 19182 17490 19234 17502
rect 20638 17554 20690 17566
rect 20638 17490 20690 17502
rect 21422 17554 21474 17566
rect 21422 17490 21474 17502
rect 22878 17554 22930 17566
rect 22878 17490 22930 17502
rect 14366 17442 14418 17454
rect 14366 17378 14418 17390
rect 21198 17442 21250 17454
rect 21198 17378 21250 17390
rect 24782 17442 24834 17454
rect 24782 17378 24834 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 15374 17106 15426 17118
rect 15374 17042 15426 17054
rect 25230 17106 25282 17118
rect 25230 17042 25282 17054
rect 25454 17106 25506 17118
rect 25454 17042 25506 17054
rect 27022 17106 27074 17118
rect 27022 17042 27074 17054
rect 15486 16994 15538 17006
rect 14130 16942 14142 16994
rect 14194 16942 14206 16994
rect 15486 16930 15538 16942
rect 26014 16994 26066 17006
rect 26014 16930 26066 16942
rect 26238 16994 26290 17006
rect 26238 16930 26290 16942
rect 26350 16994 26402 17006
rect 26350 16930 26402 16942
rect 27134 16994 27186 17006
rect 27134 16930 27186 16942
rect 25902 16882 25954 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 14914 16830 14926 16882
rect 14978 16830 14990 16882
rect 23538 16830 23550 16882
rect 23602 16830 23614 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 25902 16818 25954 16830
rect 15934 16770 15986 16782
rect 25342 16770 25394 16782
rect 12002 16718 12014 16770
rect 12066 16718 12078 16770
rect 21746 16718 21758 16770
rect 21810 16718 21822 16770
rect 15934 16706 15986 16718
rect 25342 16706 25394 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 15374 16658 15426 16670
rect 15374 16594 15426 16606
rect 40014 16658 40066 16670
rect 40014 16594 40066 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 24334 16210 24386 16222
rect 25442 16158 25454 16210
rect 25506 16158 25518 16210
rect 27570 16158 27582 16210
rect 27634 16158 27646 16210
rect 24334 16146 24386 16158
rect 14254 16098 14306 16110
rect 14254 16034 14306 16046
rect 14478 16098 14530 16110
rect 14478 16034 14530 16046
rect 14814 16098 14866 16110
rect 14814 16034 14866 16046
rect 19070 16098 19122 16110
rect 23438 16098 23490 16110
rect 23202 16046 23214 16098
rect 23266 16046 23278 16098
rect 23874 16046 23886 16098
rect 23938 16046 23950 16098
rect 24658 16046 24670 16098
rect 24722 16046 24734 16098
rect 19070 16034 19122 16046
rect 23438 16034 23490 16046
rect 18958 15986 19010 15998
rect 18958 15922 19010 15934
rect 14478 15874 14530 15886
rect 14478 15810 14530 15822
rect 18734 15874 18786 15886
rect 18734 15810 18786 15822
rect 23550 15874 23602 15886
rect 23550 15810 23602 15822
rect 23662 15874 23714 15886
rect 23662 15810 23714 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 15150 15538 15202 15550
rect 15150 15474 15202 15486
rect 17502 15538 17554 15550
rect 17502 15474 17554 15486
rect 18062 15538 18114 15550
rect 18062 15474 18114 15486
rect 18286 15426 18338 15438
rect 13906 15374 13918 15426
rect 13970 15374 13982 15426
rect 18286 15362 18338 15374
rect 19182 15426 19234 15438
rect 19182 15362 19234 15374
rect 23886 15426 23938 15438
rect 23886 15362 23938 15374
rect 19406 15314 19458 15326
rect 14690 15262 14702 15314
rect 14754 15262 14766 15314
rect 18498 15262 18510 15314
rect 18562 15262 18574 15314
rect 18722 15262 18734 15314
rect 18786 15262 18798 15314
rect 19406 15250 19458 15262
rect 19630 15314 19682 15326
rect 19630 15250 19682 15262
rect 20974 15314 21026 15326
rect 20974 15250 21026 15262
rect 21198 15314 21250 15326
rect 21646 15314 21698 15326
rect 21522 15262 21534 15314
rect 21586 15262 21598 15314
rect 21198 15250 21250 15262
rect 21646 15250 21698 15262
rect 21870 15314 21922 15326
rect 21870 15250 21922 15262
rect 17726 15202 17778 15214
rect 11778 15150 11790 15202
rect 11842 15150 11854 15202
rect 17378 15150 17390 15202
rect 17442 15150 17454 15202
rect 17726 15138 17778 15150
rect 18174 15202 18226 15214
rect 18174 15138 18226 15150
rect 19294 15202 19346 15214
rect 21746 15150 21758 15202
rect 21810 15150 21822 15202
rect 19294 15138 19346 15150
rect 23774 15090 23826 15102
rect 23774 15026 23826 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19518 14642 19570 14654
rect 16706 14590 16718 14642
rect 16770 14590 16782 14642
rect 18834 14590 18846 14642
rect 18898 14590 18910 14642
rect 19518 14578 19570 14590
rect 20526 14642 20578 14654
rect 20526 14578 20578 14590
rect 22094 14642 22146 14654
rect 23650 14590 23662 14642
rect 23714 14590 23726 14642
rect 25778 14590 25790 14642
rect 25842 14590 25854 14642
rect 22094 14578 22146 14590
rect 19294 14530 19346 14542
rect 15922 14478 15934 14530
rect 15986 14478 15998 14530
rect 19294 14466 19346 14478
rect 19966 14530 20018 14542
rect 22866 14478 22878 14530
rect 22930 14478 22942 14530
rect 19966 14466 20018 14478
rect 22430 14418 22482 14430
rect 22430 14354 22482 14366
rect 22542 14418 22594 14430
rect 22542 14354 22594 14366
rect 19742 14306 19794 14318
rect 19742 14242 19794 14254
rect 19854 14306 19906 14318
rect 19854 14242 19906 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 23998 13970 24050 13982
rect 23998 13906 24050 13918
rect 16830 13858 16882 13870
rect 18162 13806 18174 13858
rect 18226 13806 18238 13858
rect 21410 13806 21422 13858
rect 21474 13806 21486 13858
rect 16830 13794 16882 13806
rect 17378 13694 17390 13746
rect 17442 13694 17454 13746
rect 20738 13694 20750 13746
rect 20802 13694 20814 13746
rect 20290 13582 20302 13634
rect 20354 13582 20366 13634
rect 23538 13582 23550 13634
rect 23602 13582 23614 13634
rect 16718 13522 16770 13534
rect 16718 13458 16770 13470
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 20638 13186 20690 13198
rect 18610 13134 18622 13186
rect 18674 13183 18686 13186
rect 19170 13183 19182 13186
rect 18674 13137 19182 13183
rect 18674 13134 18686 13137
rect 19170 13134 19182 13137
rect 19234 13134 19246 13186
rect 20638 13122 20690 13134
rect 18622 13074 18674 13086
rect 15922 13022 15934 13074
rect 15986 13022 15998 13074
rect 18050 13022 18062 13074
rect 18114 13022 18126 13074
rect 18622 13010 18674 13022
rect 19182 13074 19234 13086
rect 19182 13010 19234 13022
rect 15138 12910 15150 12962
rect 15202 12910 15214 12962
rect 20750 12850 20802 12862
rect 20750 12786 20802 12798
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 20078 4114 20130 4126
rect 20078 4050 20130 4062
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19518 38222 19570 38274
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 14814 38110 14866 38162
rect 15934 37998 15986 38050
rect 17614 37998 17666 38050
rect 21422 37998 21474 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 21422 37438 21474 37490
rect 1710 37326 1762 37378
rect 17390 37214 17442 37266
rect 20862 37214 20914 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 16718 36654 16770 36706
rect 15710 36430 15762 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 13470 28702 13522 28754
rect 16270 28590 16322 28642
rect 16830 28590 16882 28642
rect 15598 28478 15650 28530
rect 18510 28478 18562 28530
rect 18622 28478 18674 28530
rect 18846 28366 18898 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 14926 28030 14978 28082
rect 15262 28030 15314 28082
rect 15486 28030 15538 28082
rect 15710 27918 15762 27970
rect 14142 27806 14194 27858
rect 15822 27806 15874 27858
rect 20302 27806 20354 27858
rect 11230 27694 11282 27746
rect 13358 27694 13410 27746
rect 14590 27694 14642 27746
rect 17390 27694 17442 27746
rect 19518 27694 19570 27746
rect 20750 27694 20802 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 15598 27246 15650 27298
rect 1934 27134 1986 27186
rect 4286 27022 4338 27074
rect 13918 27022 13970 27074
rect 15150 27022 15202 27074
rect 19070 27022 19122 27074
rect 19406 27022 19458 27074
rect 13806 26910 13858 26962
rect 14254 26910 14306 26962
rect 14590 26910 14642 26962
rect 14814 26910 14866 26962
rect 15038 26910 15090 26962
rect 15598 26910 15650 26962
rect 15710 26910 15762 26962
rect 21870 26910 21922 26962
rect 22094 26910 22146 26962
rect 22206 26910 22258 26962
rect 13582 26798 13634 26850
rect 14478 26798 14530 26850
rect 19182 26798 19234 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17950 26462 18002 26514
rect 13134 26350 13186 26402
rect 25566 26350 25618 26402
rect 12462 26238 12514 26290
rect 18174 26238 18226 26290
rect 20414 26238 20466 26290
rect 25342 26238 25394 26290
rect 37662 26238 37714 26290
rect 15262 26126 15314 26178
rect 15710 26126 15762 26178
rect 19518 26126 19570 26178
rect 19966 26126 20018 26178
rect 21086 26126 21138 26178
rect 23214 26126 23266 26178
rect 39902 26126 39954 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 13918 25678 13970 25730
rect 21310 25678 21362 25730
rect 21422 25678 21474 25730
rect 20638 25566 20690 25618
rect 40014 25566 40066 25618
rect 13694 25454 13746 25506
rect 17726 25454 17778 25506
rect 21870 25454 21922 25506
rect 22094 25454 22146 25506
rect 22766 25454 22818 25506
rect 37886 25454 37938 25506
rect 14254 25342 14306 25394
rect 15374 25342 15426 25394
rect 18510 25342 18562 25394
rect 21534 25342 21586 25394
rect 23550 25342 23602 25394
rect 14030 25230 14082 25282
rect 14926 25230 14978 25282
rect 15038 25230 15090 25282
rect 15150 25230 15202 25282
rect 25790 25230 25842 25282
rect 26238 25230 26290 25282
rect 26574 25230 26626 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 13470 24894 13522 24946
rect 13694 24894 13746 24946
rect 17502 24894 17554 24946
rect 23774 24894 23826 24946
rect 14702 24782 14754 24834
rect 18286 24782 18338 24834
rect 13358 24670 13410 24722
rect 14030 24670 14082 24722
rect 23326 24670 23378 24722
rect 23998 24670 24050 24722
rect 24670 24670 24722 24722
rect 25230 24670 25282 24722
rect 37662 24670 37714 24722
rect 16830 24558 16882 24610
rect 26014 24558 26066 24610
rect 28142 24558 28194 24610
rect 23662 24446 23714 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 18174 24110 18226 24162
rect 13694 23998 13746 24050
rect 19406 23998 19458 24050
rect 22430 23998 22482 24050
rect 25230 23998 25282 24050
rect 40014 23998 40066 24050
rect 13806 23886 13858 23938
rect 14366 23886 14418 23938
rect 17278 23886 17330 23938
rect 19630 23886 19682 23938
rect 20078 23886 20130 23938
rect 20190 23886 20242 23938
rect 22766 23886 22818 23938
rect 23774 23886 23826 23938
rect 23886 23886 23938 23938
rect 25118 23886 25170 23938
rect 25790 23886 25842 23938
rect 26126 23886 26178 23938
rect 37662 23886 37714 23938
rect 17838 23774 17890 23826
rect 19406 23774 19458 23826
rect 23102 23774 23154 23826
rect 23438 23774 23490 23826
rect 26350 23774 26402 23826
rect 26462 23774 26514 23826
rect 17502 23662 17554 23714
rect 18062 23662 18114 23714
rect 19966 23662 20018 23714
rect 20414 23662 20466 23714
rect 23662 23662 23714 23714
rect 25342 23662 25394 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 15374 23326 15426 23378
rect 22766 23326 22818 23378
rect 14142 23214 14194 23266
rect 14366 23214 14418 23266
rect 15150 23214 15202 23266
rect 15598 23214 15650 23266
rect 11006 23102 11058 23154
rect 14926 23102 14978 23154
rect 15710 23102 15762 23154
rect 19406 23102 19458 23154
rect 11678 22990 11730 23042
rect 13806 22990 13858 23042
rect 14254 22990 14306 23042
rect 17502 22990 17554 23042
rect 20190 22990 20242 23042
rect 22318 22990 22370 23042
rect 17614 22878 17666 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 14478 22542 14530 22594
rect 15038 22542 15090 22594
rect 15822 22542 15874 22594
rect 24894 22430 24946 22482
rect 40014 22430 40066 22482
rect 14926 22318 14978 22370
rect 16158 22318 16210 22370
rect 22766 22318 22818 22370
rect 37662 22318 37714 22370
rect 14590 22206 14642 22258
rect 15934 22206 15986 22258
rect 17390 22206 17442 22258
rect 17614 22206 17666 22258
rect 19630 22206 19682 22258
rect 19742 22206 19794 22258
rect 19966 22206 20018 22258
rect 21422 22206 21474 22258
rect 21534 22206 21586 22258
rect 22430 22206 22482 22258
rect 22542 22206 22594 22258
rect 14030 22094 14082 22146
rect 14478 22094 14530 22146
rect 17502 22094 17554 22146
rect 18174 22094 18226 22146
rect 18510 22094 18562 22146
rect 18958 22094 19010 22146
rect 20190 22094 20242 22146
rect 20526 22094 20578 22146
rect 21198 22094 21250 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14590 21758 14642 21810
rect 24334 21758 24386 21810
rect 14926 21646 14978 21698
rect 28814 21646 28866 21698
rect 4286 21534 4338 21586
rect 18622 21534 18674 21586
rect 24110 21534 24162 21586
rect 25230 21534 25282 21586
rect 28590 21534 28642 21586
rect 37662 21534 37714 21586
rect 13134 21422 13186 21474
rect 17502 21422 17554 21474
rect 17726 21422 17778 21474
rect 23438 21422 23490 21474
rect 26014 21422 26066 21474
rect 28142 21422 28194 21474
rect 40014 21422 40066 21474
rect 1934 21310 1986 21362
rect 18062 21310 18114 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 13918 20974 13970 21026
rect 15038 20974 15090 21026
rect 17950 20974 18002 21026
rect 24222 20974 24274 21026
rect 9998 20862 10050 20914
rect 17166 20862 17218 20914
rect 19966 20862 20018 20914
rect 23214 20862 23266 20914
rect 24446 20862 24498 20914
rect 24558 20862 24610 20914
rect 27022 20862 27074 20914
rect 40014 20862 40066 20914
rect 12910 20750 12962 20802
rect 13582 20750 13634 20802
rect 14478 20750 14530 20802
rect 14926 20750 14978 20802
rect 15262 20750 15314 20802
rect 16158 20750 16210 20802
rect 17390 20750 17442 20802
rect 17726 20750 17778 20802
rect 19630 20750 19682 20802
rect 20078 20750 20130 20802
rect 21310 20750 21362 20802
rect 22206 20750 22258 20802
rect 23774 20750 23826 20802
rect 37662 20750 37714 20802
rect 12126 20638 12178 20690
rect 15374 20638 15426 20690
rect 15486 20638 15538 20690
rect 15822 20638 15874 20690
rect 19854 20638 19906 20690
rect 20302 20638 20354 20690
rect 23102 20638 23154 20690
rect 23998 20638 24050 20690
rect 24670 20638 24722 20690
rect 26014 20638 26066 20690
rect 26910 20638 26962 20690
rect 13806 20526 13858 20578
rect 18846 20526 18898 20578
rect 19182 20526 19234 20578
rect 21646 20526 21698 20578
rect 21982 20526 22034 20578
rect 23326 20526 23378 20578
rect 26126 20526 26178 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14478 20190 14530 20242
rect 16382 20190 16434 20242
rect 18622 20190 18674 20242
rect 12126 20078 12178 20130
rect 14702 20078 14754 20130
rect 14814 20078 14866 20130
rect 18062 20078 18114 20130
rect 18958 20078 19010 20130
rect 20862 20078 20914 20130
rect 26238 20078 26290 20130
rect 11454 19966 11506 20018
rect 16270 19966 16322 20018
rect 18286 19966 18338 20018
rect 19742 19966 19794 20018
rect 20302 19966 20354 20018
rect 25454 19966 25506 20018
rect 14254 19854 14306 19906
rect 15374 19854 15426 19906
rect 16158 19854 16210 19906
rect 20190 19854 20242 19906
rect 21422 19854 21474 19906
rect 24782 19854 24834 19906
rect 28366 19854 28418 19906
rect 17950 19742 18002 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15822 19406 15874 19458
rect 17726 19406 17778 19458
rect 15486 19294 15538 19346
rect 16382 19294 16434 19346
rect 17838 19294 17890 19346
rect 19070 19294 19122 19346
rect 22094 19294 22146 19346
rect 24222 19294 24274 19346
rect 25454 19294 25506 19346
rect 14926 19182 14978 19234
rect 16158 19182 16210 19234
rect 17054 19182 17106 19234
rect 18062 19182 18114 19234
rect 18958 19182 19010 19234
rect 19406 19182 19458 19234
rect 21422 19182 21474 19234
rect 25118 19182 25170 19234
rect 25790 19182 25842 19234
rect 20414 19070 20466 19122
rect 25566 19070 25618 19122
rect 17390 18958 17442 19010
rect 19966 18958 20018 19010
rect 20750 18958 20802 19010
rect 25342 18958 25394 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 16830 18622 16882 18674
rect 18622 18622 18674 18674
rect 19182 18622 19234 18674
rect 22318 18622 22370 18674
rect 23550 18622 23602 18674
rect 25902 18622 25954 18674
rect 17726 18510 17778 18562
rect 18734 18510 18786 18562
rect 19070 18510 19122 18562
rect 20750 18510 20802 18562
rect 21870 18510 21922 18562
rect 22430 18510 22482 18562
rect 16494 18398 16546 18450
rect 18062 18398 18114 18450
rect 18398 18398 18450 18450
rect 19630 18398 19682 18450
rect 20078 18398 20130 18450
rect 21422 18398 21474 18450
rect 21982 18398 22034 18450
rect 23774 18398 23826 18450
rect 25230 18398 25282 18450
rect 25678 18398 25730 18450
rect 26126 18398 26178 18450
rect 37662 18398 37714 18450
rect 21310 18286 21362 18338
rect 25454 18286 25506 18338
rect 26014 18286 26066 18338
rect 21086 18174 21138 18226
rect 21870 18174 21922 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 17950 17838 18002 17890
rect 18062 17838 18114 17890
rect 18286 17838 18338 17890
rect 18846 17838 18898 17890
rect 19630 17838 19682 17890
rect 20190 17838 20242 17890
rect 20302 17838 20354 17890
rect 21982 17838 22034 17890
rect 22654 17838 22706 17890
rect 1934 17726 1986 17778
rect 15038 17726 15090 17778
rect 21870 17726 21922 17778
rect 22990 17726 23042 17778
rect 25902 17726 25954 17778
rect 28030 17726 28082 17778
rect 4286 17614 4338 17666
rect 14366 17614 14418 17666
rect 14702 17614 14754 17666
rect 15262 17614 15314 17666
rect 15486 17614 15538 17666
rect 17054 17614 17106 17666
rect 18398 17614 18450 17666
rect 19070 17614 19122 17666
rect 19406 17614 19458 17666
rect 20526 17614 20578 17666
rect 21534 17614 21586 17666
rect 25118 17614 25170 17666
rect 14030 17502 14082 17554
rect 14926 17502 14978 17554
rect 17390 17502 17442 17554
rect 19182 17502 19234 17554
rect 20638 17502 20690 17554
rect 21422 17502 21474 17554
rect 22878 17502 22930 17554
rect 14366 17390 14418 17442
rect 21198 17390 21250 17442
rect 24782 17390 24834 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 15374 17054 15426 17106
rect 25230 17054 25282 17106
rect 25454 17054 25506 17106
rect 27022 17054 27074 17106
rect 14142 16942 14194 16994
rect 15486 16942 15538 16994
rect 26014 16942 26066 16994
rect 26238 16942 26290 16994
rect 26350 16942 26402 16994
rect 27134 16942 27186 16994
rect 4286 16830 4338 16882
rect 14926 16830 14978 16882
rect 23550 16830 23602 16882
rect 25902 16830 25954 16882
rect 37662 16830 37714 16882
rect 12014 16718 12066 16770
rect 15934 16718 15986 16770
rect 21758 16718 21810 16770
rect 25342 16718 25394 16770
rect 1934 16606 1986 16658
rect 15374 16606 15426 16658
rect 40014 16606 40066 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 24334 16158 24386 16210
rect 25454 16158 25506 16210
rect 27582 16158 27634 16210
rect 14254 16046 14306 16098
rect 14478 16046 14530 16098
rect 14814 16046 14866 16098
rect 19070 16046 19122 16098
rect 23214 16046 23266 16098
rect 23438 16046 23490 16098
rect 23886 16046 23938 16098
rect 24670 16046 24722 16098
rect 18958 15934 19010 15986
rect 14478 15822 14530 15874
rect 18734 15822 18786 15874
rect 23550 15822 23602 15874
rect 23662 15822 23714 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 15150 15486 15202 15538
rect 17502 15486 17554 15538
rect 18062 15486 18114 15538
rect 13918 15374 13970 15426
rect 18286 15374 18338 15426
rect 19182 15374 19234 15426
rect 23886 15374 23938 15426
rect 14702 15262 14754 15314
rect 18510 15262 18562 15314
rect 18734 15262 18786 15314
rect 19406 15262 19458 15314
rect 19630 15262 19682 15314
rect 20974 15262 21026 15314
rect 21198 15262 21250 15314
rect 21534 15262 21586 15314
rect 21646 15262 21698 15314
rect 21870 15262 21922 15314
rect 11790 15150 11842 15202
rect 17390 15150 17442 15202
rect 17726 15150 17778 15202
rect 18174 15150 18226 15202
rect 19294 15150 19346 15202
rect 21758 15150 21810 15202
rect 23774 15038 23826 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 16718 14590 16770 14642
rect 18846 14590 18898 14642
rect 19518 14590 19570 14642
rect 20526 14590 20578 14642
rect 22094 14590 22146 14642
rect 23662 14590 23714 14642
rect 25790 14590 25842 14642
rect 15934 14478 15986 14530
rect 19294 14478 19346 14530
rect 19966 14478 20018 14530
rect 22878 14478 22930 14530
rect 22430 14366 22482 14418
rect 22542 14366 22594 14418
rect 19742 14254 19794 14306
rect 19854 14254 19906 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 23998 13918 24050 13970
rect 16830 13806 16882 13858
rect 18174 13806 18226 13858
rect 21422 13806 21474 13858
rect 17390 13694 17442 13746
rect 20750 13694 20802 13746
rect 20302 13582 20354 13634
rect 23550 13582 23602 13634
rect 16718 13470 16770 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 18622 13134 18674 13186
rect 19182 13134 19234 13186
rect 20638 13134 20690 13186
rect 15934 13022 15986 13074
rect 18062 13022 18114 13074
rect 18622 13022 18674 13074
rect 19182 13022 19234 13074
rect 15150 12910 15202 12962
rect 20750 12798 20802 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 19070 4286 19122 4338
rect 25230 4286 25282 4338
rect 20078 4062 20130 4114
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 22094 3614 22146 3666
rect 25566 3614 25618 3666
rect 17614 3502 17666 3554
rect 21086 3502 21138 3554
rect 24558 3502 24610 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 14784 41200 14896 42000
rect 15456 41200 15568 42000
rect 16128 41200 16240 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 14812 38162 14868 41200
rect 14812 38110 14814 38162
rect 14866 38110 14868 38162
rect 14812 38098 14868 38110
rect 14924 38052 14980 38062
rect 1708 37378 1764 37390
rect 1708 37326 1710 37378
rect 1762 37326 1764 37378
rect 1708 37044 1764 37326
rect 1708 36978 1764 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 13468 28754 13524 28766
rect 13468 28702 13470 28754
rect 13522 28702 13524 28754
rect 13468 28532 13524 28702
rect 13468 28466 13524 28476
rect 14588 28644 14644 28654
rect 4172 28308 4228 28318
rect 1932 27188 1988 27198
rect 1932 27094 1988 27132
rect 4172 22148 4228 28252
rect 14140 27858 14196 27870
rect 14140 27806 14142 27858
rect 14194 27806 14196 27858
rect 11228 27746 11284 27758
rect 11228 27694 11230 27746
rect 11282 27694 11284 27746
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 11228 27076 11284 27694
rect 11228 27010 11284 27020
rect 13356 27746 13412 27758
rect 13356 27694 13358 27746
rect 13410 27694 13412 27746
rect 13132 26964 13188 26974
rect 13132 26402 13188 26908
rect 13132 26350 13134 26402
rect 13186 26350 13188 26402
rect 13132 26338 13188 26350
rect 12460 26290 12516 26302
rect 12460 26238 12462 26290
rect 12514 26238 12516 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 12460 25284 12516 26238
rect 13356 25732 13412 27694
rect 14140 27748 14196 27806
rect 14588 27748 14644 28588
rect 14140 27746 14644 27748
rect 14140 27694 14590 27746
rect 14642 27694 14644 27746
rect 14140 27692 14644 27694
rect 13916 27188 13972 27198
rect 13804 27076 13860 27086
rect 13804 26962 13860 27020
rect 13916 27074 13972 27132
rect 13916 27022 13918 27074
rect 13970 27022 13972 27074
rect 13916 27010 13972 27022
rect 13804 26910 13806 26962
rect 13858 26910 13860 26962
rect 13804 26898 13860 26910
rect 13356 25666 13412 25676
rect 13580 26850 13636 26862
rect 13580 26798 13582 26850
rect 13634 26798 13636 26850
rect 13580 25508 13636 26798
rect 14140 26180 14196 27692
rect 14588 27682 14644 27692
rect 14924 28532 14980 37996
rect 15484 36708 15540 41200
rect 15932 38052 15988 38062
rect 15932 37958 15988 37996
rect 16156 37492 16212 41200
rect 19516 38274 19572 41200
rect 19516 38222 19518 38274
rect 19570 38222 19572 38274
rect 19516 38210 19572 38222
rect 16156 37426 16212 37436
rect 17612 38050 17668 38062
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 17388 37268 17444 37278
rect 17276 37266 17444 37268
rect 17276 37214 17390 37266
rect 17442 37214 17444 37266
rect 17276 37212 17444 37214
rect 15484 36642 15540 36652
rect 16716 36708 16772 36718
rect 16716 36614 16772 36652
rect 15708 36482 15764 36494
rect 15708 36430 15710 36482
rect 15762 36430 15764 36482
rect 15708 31948 15764 36430
rect 14924 28082 14980 28476
rect 14924 28030 14926 28082
rect 14978 28030 14980 28082
rect 14364 27524 14420 27534
rect 14252 26964 14308 26974
rect 14252 26870 14308 26908
rect 13916 25732 13972 25742
rect 13916 25638 13972 25676
rect 13692 25508 13748 25518
rect 13580 25506 13748 25508
rect 13580 25454 13694 25506
rect 13746 25454 13748 25506
rect 13580 25452 13748 25454
rect 13692 25442 13748 25452
rect 14028 25284 14084 25294
rect 12460 25218 12516 25228
rect 13692 25282 14084 25284
rect 13692 25230 14030 25282
rect 14082 25230 14084 25282
rect 13692 25228 14084 25230
rect 13468 24948 13524 24958
rect 13468 24854 13524 24892
rect 13692 24946 13748 25228
rect 14028 25218 14084 25228
rect 13692 24894 13694 24946
rect 13746 24894 13748 24946
rect 13692 24882 13748 24894
rect 14028 25060 14084 25070
rect 14140 25060 14196 26124
rect 14252 25396 14308 25406
rect 14364 25396 14420 27468
rect 14924 27076 14980 28030
rect 15260 31892 15764 31948
rect 15260 28082 15316 31892
rect 16268 28644 16324 28654
rect 16268 28550 16324 28588
rect 16828 28644 16884 28654
rect 16828 28550 16884 28588
rect 15596 28530 15652 28542
rect 15596 28478 15598 28530
rect 15650 28478 15652 28530
rect 15260 28030 15262 28082
rect 15314 28030 15316 28082
rect 15260 28018 15316 28030
rect 15484 28084 15540 28094
rect 15596 28084 15652 28478
rect 15484 28082 15652 28084
rect 15484 28030 15486 28082
rect 15538 28030 15652 28082
rect 15484 28028 15652 28030
rect 15484 28018 15540 28028
rect 15708 27970 15764 27982
rect 15708 27918 15710 27970
rect 15762 27918 15764 27970
rect 15708 27524 15764 27918
rect 15708 27458 15764 27468
rect 15820 27858 15876 27870
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 15596 27300 15652 27310
rect 15820 27300 15876 27806
rect 15596 27298 15876 27300
rect 15596 27246 15598 27298
rect 15650 27246 15876 27298
rect 15596 27244 15876 27246
rect 15596 27234 15652 27244
rect 14924 27010 14980 27020
rect 15148 27188 15204 27198
rect 15148 27074 15204 27132
rect 15148 27022 15150 27074
rect 15202 27022 15204 27074
rect 15148 27010 15204 27022
rect 15596 27076 15652 27086
rect 15820 27076 15876 27086
rect 14588 26964 14644 26974
rect 14812 26964 14868 26974
rect 14588 26962 14868 26964
rect 14588 26910 14590 26962
rect 14642 26910 14814 26962
rect 14866 26910 14868 26962
rect 14588 26908 14868 26910
rect 14588 26898 14644 26908
rect 14812 26898 14868 26908
rect 15036 26964 15092 26974
rect 14476 26852 14532 26862
rect 14476 26758 14532 26796
rect 15036 26740 15092 26908
rect 15596 26962 15652 27020
rect 15596 26910 15598 26962
rect 15650 26910 15652 26962
rect 15596 26898 15652 26910
rect 15708 27020 15820 27076
rect 15708 26962 15764 27020
rect 15820 27010 15876 27020
rect 15708 26910 15710 26962
rect 15762 26910 15764 26962
rect 15708 26898 15764 26910
rect 17276 26964 17332 37212
rect 17388 37202 17444 37212
rect 17612 31948 17668 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 20188 37492 20244 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 22876 38276 22932 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 22876 38210 22932 38220
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 21420 38052 21476 38062
rect 20188 37426 20244 37436
rect 20972 38050 21476 38052
rect 20972 37998 21422 38050
rect 21474 37998 21476 38050
rect 20972 37996 21476 37998
rect 20860 37266 20916 37278
rect 20860 37214 20862 37266
rect 20914 37214 20916 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 17388 31892 17668 31948
rect 17388 28532 17444 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 18508 28532 18564 28542
rect 17388 27746 17444 28476
rect 17388 27694 17390 27746
rect 17442 27694 17444 27746
rect 17388 27682 17444 27694
rect 17948 28530 18564 28532
rect 17948 28478 18510 28530
rect 18562 28478 18564 28530
rect 17948 28476 18564 28478
rect 17276 26898 17332 26908
rect 17948 27076 18004 28476
rect 18508 28466 18564 28476
rect 18620 28532 18676 28542
rect 18620 28438 18676 28476
rect 18844 28420 18900 28430
rect 18844 28418 19124 28420
rect 18844 28366 18846 28418
rect 18898 28366 19124 28418
rect 18844 28364 19124 28366
rect 18844 28354 18900 28364
rect 15372 26852 15428 26862
rect 15036 26684 15316 26740
rect 15260 26178 15316 26684
rect 15260 26126 15262 26178
rect 15314 26126 15316 26178
rect 15260 26114 15316 26126
rect 14252 25394 14532 25396
rect 14252 25342 14254 25394
rect 14306 25342 14532 25394
rect 14252 25340 14532 25342
rect 14252 25330 14308 25340
rect 14084 25004 14196 25060
rect 13356 24722 13412 24734
rect 13356 24670 13358 24722
rect 13410 24670 13412 24722
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 13356 24164 13412 24670
rect 14028 24722 14084 25004
rect 14028 24670 14030 24722
rect 14082 24670 14084 24722
rect 13356 24108 13748 24164
rect 13692 24050 13748 24108
rect 13692 23998 13694 24050
rect 13746 23998 13748 24050
rect 13692 23716 13748 23998
rect 13692 23650 13748 23660
rect 13804 23940 13860 23950
rect 13804 23268 13860 23884
rect 13692 23212 13860 23268
rect 11004 23154 11060 23166
rect 11004 23102 11006 23154
rect 11058 23102 11060 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 22082 4228 22092
rect 11004 22036 11060 23102
rect 11676 23044 11732 23054
rect 11676 22950 11732 22988
rect 11004 21970 11060 21980
rect 13132 22036 13188 22046
rect 4284 21588 4340 21598
rect 4284 21494 4340 21532
rect 9996 21588 10052 21598
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1932 20850 1988 20860
rect 9996 20916 10052 21532
rect 9996 20822 10052 20860
rect 13132 21474 13188 21980
rect 13132 21422 13134 21474
rect 13186 21422 13188 21474
rect 12908 20804 12964 20814
rect 13132 20804 13188 21422
rect 12908 20802 13188 20804
rect 12908 20750 12910 20802
rect 12962 20750 13188 20802
rect 12908 20748 13188 20750
rect 13580 20804 13636 20814
rect 13692 20804 13748 23212
rect 13804 23042 13860 23054
rect 13804 22990 13806 23042
rect 13858 22990 13860 23042
rect 13804 22932 13860 22990
rect 13916 22932 13972 22942
rect 13804 22876 13916 22932
rect 13916 22866 13972 22876
rect 14028 22146 14084 24670
rect 14364 23938 14420 23950
rect 14364 23886 14366 23938
rect 14418 23886 14420 23938
rect 14364 23828 14420 23886
rect 14364 23762 14420 23772
rect 14140 23716 14196 23726
rect 14140 23266 14196 23660
rect 14140 23214 14142 23266
rect 14194 23214 14196 23266
rect 14140 23202 14196 23214
rect 14364 23266 14420 23278
rect 14364 23214 14366 23266
rect 14418 23214 14420 23266
rect 14252 23044 14308 23054
rect 14252 22950 14308 22988
rect 14028 22094 14030 22146
rect 14082 22094 14084 22146
rect 14028 22036 14084 22094
rect 14028 21970 14084 21980
rect 13916 21924 13972 21934
rect 13916 21026 13972 21868
rect 13916 20974 13918 21026
rect 13970 20974 13972 21026
rect 13916 20962 13972 20974
rect 14028 21700 14084 21710
rect 14364 21700 14420 23214
rect 14476 22594 14532 25340
rect 15372 25394 15428 26796
rect 17948 26514 18004 27020
rect 19068 27074 19124 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20300 27858 20356 27870
rect 20300 27806 20302 27858
rect 20354 27806 20356 27858
rect 19516 27748 19572 27758
rect 19068 27022 19070 27074
rect 19122 27022 19124 27074
rect 19068 27010 19124 27022
rect 19404 27746 19572 27748
rect 19404 27694 19518 27746
rect 19570 27694 19572 27746
rect 19404 27692 19572 27694
rect 19404 27074 19460 27692
rect 19516 27682 19572 27692
rect 20300 27748 20356 27806
rect 20748 27748 20804 27758
rect 20300 27746 20804 27748
rect 20300 27694 20750 27746
rect 20802 27694 20804 27746
rect 20300 27692 20804 27694
rect 19404 27022 19406 27074
rect 19458 27022 19460 27074
rect 19404 27010 19460 27022
rect 20300 26908 20356 27692
rect 20748 27682 20804 27692
rect 20860 26908 20916 37214
rect 19180 26852 19236 26862
rect 20300 26852 20468 26908
rect 19180 26850 19460 26852
rect 19180 26798 19182 26850
rect 19234 26798 19460 26850
rect 19180 26796 19460 26798
rect 19180 26786 19236 26796
rect 17948 26462 17950 26514
rect 18002 26462 18004 26514
rect 17948 26450 18004 26462
rect 18172 26290 18228 26302
rect 18172 26238 18174 26290
rect 18226 26238 18228 26290
rect 15708 26180 15764 26190
rect 15708 26086 15764 26124
rect 17724 26180 17780 26190
rect 17724 25508 17780 26124
rect 15372 25342 15374 25394
rect 15426 25342 15428 25394
rect 14924 25282 14980 25294
rect 14924 25230 14926 25282
rect 14978 25230 14980 25282
rect 14924 25060 14980 25230
rect 14588 25004 14980 25060
rect 15036 25282 15092 25294
rect 15036 25230 15038 25282
rect 15090 25230 15092 25282
rect 14588 23940 14644 25004
rect 15036 24948 15092 25230
rect 14700 24892 15092 24948
rect 15148 25282 15204 25294
rect 15148 25230 15150 25282
rect 15202 25230 15204 25282
rect 15148 24948 15204 25230
rect 14700 24834 14756 24892
rect 14700 24782 14702 24834
rect 14754 24782 14756 24834
rect 14700 24770 14756 24782
rect 14588 23874 14644 23884
rect 15036 23828 15092 23838
rect 14476 22542 14478 22594
rect 14530 22542 14532 22594
rect 14476 22530 14532 22542
rect 14924 23154 14980 23166
rect 14924 23102 14926 23154
rect 14978 23102 14980 23154
rect 14924 22932 14980 23102
rect 14924 22370 14980 22876
rect 14924 22318 14926 22370
rect 14978 22318 14980 22370
rect 14924 22306 14980 22318
rect 15036 22594 15092 23772
rect 15148 23716 15204 24892
rect 15148 23650 15204 23660
rect 15372 23378 15428 25342
rect 17500 25506 17780 25508
rect 17500 25454 17726 25506
rect 17778 25454 17780 25506
rect 17500 25452 17780 25454
rect 17500 24946 17556 25452
rect 17724 25442 17780 25452
rect 17500 24894 17502 24946
rect 17554 24894 17556 24946
rect 17500 24836 17556 24894
rect 17500 24770 17556 24780
rect 18172 24948 18228 26238
rect 19404 25508 19460 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20412 26290 20468 26852
rect 20412 26238 20414 26290
rect 20466 26238 20468 26290
rect 19516 26180 19572 26190
rect 19516 26086 19572 26124
rect 19964 26180 20020 26190
rect 19964 26086 20020 26124
rect 20412 26180 20468 26238
rect 20412 26114 20468 26124
rect 20636 26852 20916 26908
rect 20636 25618 20692 26852
rect 20636 25566 20638 25618
rect 20690 25566 20692 25618
rect 19404 25452 19572 25508
rect 18508 25396 18564 25406
rect 18508 25394 19460 25396
rect 18508 25342 18510 25394
rect 18562 25342 19460 25394
rect 18508 25340 19460 25342
rect 18508 25330 18564 25340
rect 16828 24612 16884 24622
rect 16828 24610 17220 24612
rect 16828 24558 16830 24610
rect 16882 24558 17220 24610
rect 16828 24556 17220 24558
rect 16828 24546 16884 24556
rect 15372 23326 15374 23378
rect 15426 23326 15428 23378
rect 15372 23314 15428 23326
rect 15148 23268 15204 23278
rect 15148 23174 15204 23212
rect 15596 23266 15652 23278
rect 15596 23214 15598 23266
rect 15650 23214 15652 23266
rect 15036 22542 15038 22594
rect 15090 22542 15092 22594
rect 14588 22260 14644 22270
rect 14476 22146 14532 22158
rect 14476 22094 14478 22146
rect 14530 22094 14532 22146
rect 14476 22036 14532 22094
rect 14476 21970 14532 21980
rect 14588 21812 14644 22204
rect 14588 21810 14868 21812
rect 14588 21758 14590 21810
rect 14642 21758 14868 21810
rect 14588 21756 14868 21758
rect 14588 21746 14644 21756
rect 14476 21700 14532 21710
rect 14364 21644 14476 21700
rect 13636 20748 13748 20804
rect 12908 20738 12964 20748
rect 13580 20710 13636 20748
rect 12124 20692 12180 20702
rect 12124 20598 12180 20636
rect 12236 20580 12292 20590
rect 12236 20188 12292 20524
rect 13804 20580 13860 20590
rect 13804 20486 13860 20524
rect 12124 20132 12292 20188
rect 12124 20130 12180 20132
rect 12124 20078 12126 20130
rect 12178 20078 12180 20130
rect 12124 20066 12180 20078
rect 11452 20018 11508 20030
rect 11452 19966 11454 20018
rect 11506 19966 11508 20018
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 11452 18452 11508 19966
rect 11452 18386 11508 18396
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17778 1988 17790
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 16884 1988 17726
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 12012 17668 12068 17678
rect 1932 16818 1988 16828
rect 4284 16996 4340 17006
rect 4284 16882 4340 16940
rect 4284 16830 4286 16882
rect 4338 16830 4340 16882
rect 4284 16818 4340 16830
rect 11788 16996 11844 17006
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1932 16146 1988 16156
rect 11788 15202 11844 16940
rect 12012 16770 12068 17612
rect 12012 16718 12014 16770
rect 12066 16718 12068 16770
rect 12012 16706 12068 16718
rect 14028 17554 14084 21644
rect 14476 21634 14532 21644
rect 14812 21476 14868 21756
rect 14924 21700 14980 21710
rect 14924 21606 14980 21644
rect 15036 21588 15092 22542
rect 15036 21532 15204 21588
rect 14812 21420 15092 21476
rect 15036 21026 15092 21420
rect 15036 20974 15038 21026
rect 15090 20974 15092 21026
rect 15036 20962 15092 20974
rect 14700 20916 14756 20926
rect 14476 20802 14532 20814
rect 14476 20750 14478 20802
rect 14530 20750 14532 20802
rect 14476 20242 14532 20750
rect 14476 20190 14478 20242
rect 14530 20190 14532 20242
rect 14476 20178 14532 20190
rect 14700 20130 14756 20860
rect 14924 20802 14980 20814
rect 15148 20804 15204 21532
rect 15596 21252 15652 23214
rect 15820 23268 15876 23278
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 14700 20078 14702 20130
rect 14754 20078 14756 20130
rect 14700 20066 14756 20078
rect 14812 20468 14868 20478
rect 14812 20130 14868 20412
rect 14812 20078 14814 20130
rect 14866 20078 14868 20130
rect 14812 20066 14868 20078
rect 14252 19906 14308 19918
rect 14252 19854 14254 19906
rect 14306 19854 14308 19906
rect 14252 19236 14308 19854
rect 14252 19170 14308 19180
rect 14364 19460 14420 19470
rect 14364 17666 14420 19404
rect 14924 19460 14980 20750
rect 14924 19394 14980 19404
rect 15036 20748 15204 20804
rect 15260 21196 15652 21252
rect 15708 23154 15764 23166
rect 15708 23102 15710 23154
rect 15762 23102 15764 23154
rect 15260 20802 15316 21196
rect 15260 20750 15262 20802
rect 15314 20750 15316 20802
rect 14924 19236 14980 19246
rect 14924 19142 14980 19180
rect 15036 18788 15092 20748
rect 15260 20132 15316 20750
rect 15708 20804 15764 23102
rect 15820 22594 15876 23212
rect 17164 23044 17220 24556
rect 18172 24162 18228 24892
rect 18284 24836 18340 24846
rect 18284 24742 18340 24780
rect 19292 24836 19348 24846
rect 18172 24110 18174 24162
rect 18226 24110 18228 24162
rect 18172 24098 18228 24110
rect 17276 23940 17332 23950
rect 17276 23938 17668 23940
rect 17276 23886 17278 23938
rect 17330 23886 17668 23938
rect 17276 23884 17668 23886
rect 17276 23874 17332 23884
rect 17500 23716 17556 23726
rect 17500 23622 17556 23660
rect 17612 23492 17668 23884
rect 17836 23828 17892 23838
rect 17836 23734 17892 23772
rect 18060 23714 18116 23726
rect 18060 23662 18062 23714
rect 18114 23662 18116 23714
rect 18060 23492 18116 23662
rect 17612 23436 18116 23492
rect 17500 23044 17556 23054
rect 17164 22988 17500 23044
rect 17500 22950 17556 22988
rect 15820 22542 15822 22594
rect 15874 22542 15876 22594
rect 15820 21924 15876 22542
rect 17612 22930 17668 23436
rect 19292 23156 19348 24780
rect 19404 24050 19460 25340
rect 19404 23998 19406 24050
rect 19458 23998 19460 24050
rect 19404 23986 19460 23998
rect 19404 23828 19460 23838
rect 19404 23734 19460 23772
rect 19404 23156 19460 23166
rect 19292 23154 19460 23156
rect 19292 23102 19406 23154
rect 19458 23102 19460 23154
rect 19292 23100 19460 23102
rect 19404 23090 19460 23100
rect 17612 22878 17614 22930
rect 17666 22878 17668 22930
rect 16156 22372 16212 22382
rect 16156 22278 16212 22316
rect 17612 22372 17668 22878
rect 15932 22260 15988 22270
rect 15932 22166 15988 22204
rect 17164 22260 17220 22270
rect 15820 21858 15876 21868
rect 17164 22036 17220 22204
rect 17388 22260 17444 22270
rect 17388 22166 17444 22204
rect 17612 22258 17668 22316
rect 17612 22206 17614 22258
rect 17666 22206 17668 22258
rect 17612 22194 17668 22206
rect 18172 23044 18228 23054
rect 16380 20916 16436 20926
rect 16156 20804 16212 20814
rect 15372 20692 15428 20702
rect 15372 20598 15428 20636
rect 15484 20690 15540 20702
rect 15484 20638 15486 20690
rect 15538 20638 15540 20690
rect 15260 20066 15316 20076
rect 14924 18732 15092 18788
rect 15372 19906 15428 19918
rect 15372 19854 15374 19906
rect 15426 19854 15428 19906
rect 14924 18340 14980 18732
rect 15036 18452 15092 18462
rect 15372 18452 15428 19854
rect 15484 19460 15540 20638
rect 15708 20692 15764 20748
rect 15932 20748 16156 20804
rect 15820 20692 15876 20702
rect 15708 20690 15876 20692
rect 15708 20638 15822 20690
rect 15874 20638 15876 20690
rect 15708 20636 15876 20638
rect 15820 20626 15876 20636
rect 15484 19346 15540 19404
rect 15820 19460 15876 19470
rect 15932 19460 15988 20748
rect 16156 20710 16212 20748
rect 16380 20242 16436 20860
rect 17164 20916 17220 21980
rect 17500 22146 17556 22158
rect 17500 22094 17502 22146
rect 17554 22094 17556 22146
rect 17500 22036 17556 22094
rect 17500 21970 17556 21980
rect 18172 22146 18228 22988
rect 18172 22094 18174 22146
rect 18226 22094 18228 22146
rect 17500 21474 17556 21486
rect 17500 21422 17502 21474
rect 17554 21422 17556 21474
rect 17500 21364 17556 21422
rect 17724 21476 17780 21486
rect 17724 21382 17780 21420
rect 17500 21298 17556 21308
rect 18060 21362 18116 21374
rect 18060 21310 18062 21362
rect 18114 21310 18116 21362
rect 17948 21028 18004 21038
rect 17164 20822 17220 20860
rect 17612 20972 17948 21028
rect 17388 20804 17444 20814
rect 17388 20710 17444 20748
rect 16380 20190 16382 20242
rect 16434 20190 16436 20242
rect 16380 20178 16436 20190
rect 16268 20018 16324 20030
rect 16268 19966 16270 20018
rect 16322 19966 16324 20018
rect 15820 19458 15988 19460
rect 15820 19406 15822 19458
rect 15874 19406 15988 19458
rect 15820 19404 15988 19406
rect 16156 19906 16212 19918
rect 16156 19854 16158 19906
rect 16210 19854 16212 19906
rect 15820 19394 15876 19404
rect 15484 19294 15486 19346
rect 15538 19294 15540 19346
rect 15484 19282 15540 19294
rect 16156 19236 16212 19854
rect 16268 19348 16324 19966
rect 17612 19460 17668 20972
rect 17948 20934 18004 20972
rect 17724 20804 17780 20814
rect 18060 20804 18116 21310
rect 18172 21364 18228 22094
rect 18172 21298 18228 21308
rect 18508 22260 18564 22270
rect 18508 22146 18564 22204
rect 18508 22094 18510 22146
rect 18562 22094 18564 22146
rect 17724 20802 18116 20804
rect 17724 20750 17726 20802
rect 17778 20750 18116 20802
rect 17724 20748 18116 20750
rect 18508 20804 18564 22094
rect 18620 22148 18676 22158
rect 18956 22148 19012 22158
rect 18676 22146 19012 22148
rect 18676 22094 18958 22146
rect 19010 22094 19012 22146
rect 18676 22092 19012 22094
rect 18620 21586 18676 22092
rect 18956 22082 19012 22092
rect 19292 22036 19348 22046
rect 19348 21980 19460 22036
rect 19292 21970 19348 21980
rect 18620 21534 18622 21586
rect 18674 21534 18676 21586
rect 18620 21522 18676 21534
rect 17724 20244 17780 20748
rect 17724 20178 17780 20188
rect 18060 20132 18116 20142
rect 18060 20038 18116 20076
rect 18284 20018 18340 20030
rect 18284 19966 18286 20018
rect 18338 19966 18340 20018
rect 18284 19908 18340 19966
rect 18508 19908 18564 20748
rect 18620 21364 18676 21374
rect 18620 20242 18676 21308
rect 18620 20190 18622 20242
rect 18674 20190 18676 20242
rect 18620 20178 18676 20190
rect 18732 20692 18788 20702
rect 18284 19852 18564 19908
rect 17948 19796 18004 19806
rect 17948 19794 18340 19796
rect 17948 19742 17950 19794
rect 18002 19742 18340 19794
rect 17948 19740 18340 19742
rect 17948 19730 18004 19740
rect 17724 19460 17780 19470
rect 17612 19458 17780 19460
rect 17612 19406 17726 19458
rect 17778 19406 17780 19458
rect 17612 19404 17780 19406
rect 17724 19394 17780 19404
rect 16380 19348 16436 19358
rect 16268 19346 16436 19348
rect 16268 19294 16382 19346
rect 16434 19294 16436 19346
rect 16268 19292 16436 19294
rect 16156 19142 16212 19180
rect 16380 19124 16436 19292
rect 17836 19348 17892 19358
rect 17836 19254 17892 19292
rect 17052 19236 17108 19246
rect 17052 19142 17108 19180
rect 18060 19236 18116 19246
rect 18060 19142 18116 19180
rect 16380 19058 16436 19068
rect 17388 19010 17444 19022
rect 17388 18958 17390 19010
rect 17442 18958 17444 19010
rect 17388 18900 17444 18958
rect 17388 18834 17444 18844
rect 18060 19012 18116 19022
rect 16828 18788 16884 18798
rect 16828 18674 16884 18732
rect 16828 18622 16830 18674
rect 16882 18622 16884 18674
rect 16828 18610 16884 18622
rect 17724 18562 17780 18574
rect 17724 18510 17726 18562
rect 17778 18510 17780 18562
rect 15092 18396 15428 18452
rect 16492 18450 16548 18462
rect 16492 18398 16494 18450
rect 16546 18398 16548 18450
rect 15036 18386 15092 18396
rect 14924 18274 14980 18284
rect 15036 17780 15092 17790
rect 14364 17614 14366 17666
rect 14418 17614 14420 17666
rect 14364 17602 14420 17614
rect 14700 17778 15092 17780
rect 14700 17726 15038 17778
rect 15090 17726 15092 17778
rect 14700 17724 15092 17726
rect 14700 17666 14756 17724
rect 15036 17714 15092 17724
rect 14700 17614 14702 17666
rect 14754 17614 14756 17666
rect 14700 17602 14756 17614
rect 14028 17502 14030 17554
rect 14082 17502 14084 17554
rect 14028 16100 14084 17502
rect 14924 17554 14980 17566
rect 14924 17502 14926 17554
rect 14978 17502 14980 17554
rect 14364 17442 14420 17454
rect 14364 17390 14366 17442
rect 14418 17390 14420 17442
rect 14364 17108 14420 17390
rect 14924 17444 14980 17502
rect 14924 17378 14980 17388
rect 14140 17052 14420 17108
rect 14140 16994 14196 17052
rect 14140 16942 14142 16994
rect 14194 16942 14196 16994
rect 14140 16930 14196 16942
rect 14812 16996 14868 17006
rect 14476 16884 14532 16894
rect 14252 16100 14308 16110
rect 14028 16044 14252 16100
rect 14252 16006 14308 16044
rect 14476 16098 14532 16828
rect 14476 16046 14478 16098
rect 14530 16046 14532 16098
rect 14476 16034 14532 16046
rect 14812 16098 14868 16940
rect 14924 16884 14980 16894
rect 15148 16884 15204 18396
rect 16492 18340 16548 18398
rect 16492 18274 16548 18284
rect 17052 18340 17108 18350
rect 15484 17892 15540 17902
rect 15260 17668 15316 17678
rect 15260 17574 15316 17612
rect 15484 17666 15540 17836
rect 15484 17614 15486 17666
rect 15538 17614 15540 17666
rect 15484 17602 15540 17614
rect 17052 17666 17108 18284
rect 17724 18340 17780 18510
rect 17052 17614 17054 17666
rect 17106 17614 17108 17666
rect 17052 17602 17108 17614
rect 17388 17668 17444 17678
rect 17388 17556 17444 17612
rect 17388 17554 17556 17556
rect 17388 17502 17390 17554
rect 17442 17502 17556 17554
rect 17388 17500 17556 17502
rect 17388 17490 17444 17500
rect 15484 17444 15540 17454
rect 15372 17108 15428 17118
rect 15372 17014 15428 17052
rect 15484 16994 15540 17388
rect 15484 16942 15486 16994
rect 15538 16942 15540 16994
rect 15484 16930 15540 16942
rect 14924 16882 15204 16884
rect 14924 16830 14926 16882
rect 14978 16830 15204 16882
rect 14924 16828 15204 16830
rect 14924 16818 14980 16828
rect 14812 16046 14814 16098
rect 14866 16046 14868 16098
rect 14812 16034 14868 16046
rect 15148 16772 15204 16828
rect 14476 15874 14532 15886
rect 14476 15822 14478 15874
rect 14530 15822 14532 15874
rect 14476 15540 14532 15822
rect 15148 15540 15204 16716
rect 15372 16884 15428 16894
rect 15372 16658 15428 16828
rect 15372 16606 15374 16658
rect 15426 16606 15428 16658
rect 15372 16594 15428 16606
rect 15932 16772 15988 16782
rect 13916 15484 14532 15540
rect 14700 15538 15204 15540
rect 14700 15486 15150 15538
rect 15202 15486 15204 15538
rect 14700 15484 15204 15486
rect 13916 15426 13972 15484
rect 13916 15374 13918 15426
rect 13970 15374 13972 15426
rect 13916 15362 13972 15374
rect 14700 15314 14756 15484
rect 14700 15262 14702 15314
rect 14754 15262 14756 15314
rect 14700 15250 14756 15262
rect 11788 15150 11790 15202
rect 11842 15150 11844 15202
rect 11788 15138 11844 15150
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 15148 12962 15204 15484
rect 15932 14532 15988 16716
rect 17500 15540 17556 17500
rect 17724 17444 17780 18284
rect 17948 18452 18004 18462
rect 17948 17892 18004 18396
rect 17948 17798 18004 17836
rect 18060 18450 18116 18956
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 18060 17890 18116 18398
rect 18060 17838 18062 17890
rect 18114 17838 18116 17890
rect 18060 17826 18116 17838
rect 18284 18788 18340 19740
rect 18284 17890 18340 18732
rect 18508 18564 18564 19852
rect 18732 19348 18788 20636
rect 18844 20578 18900 20590
rect 18844 20526 18846 20578
rect 18898 20526 18900 20578
rect 18844 20244 18900 20526
rect 19180 20578 19236 20590
rect 19180 20526 19182 20578
rect 19234 20526 19236 20578
rect 19180 20468 19236 20526
rect 19180 20402 19236 20412
rect 18844 20178 18900 20188
rect 18620 19292 18788 19348
rect 18956 20130 19012 20142
rect 18956 20078 18958 20130
rect 19010 20078 19012 20130
rect 18956 20020 19012 20078
rect 18620 18674 18676 19292
rect 18956 19234 19012 19964
rect 19404 19460 19460 21980
rect 19516 20804 19572 25452
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 23940 19684 23950
rect 20076 23940 20132 23950
rect 19628 23938 20132 23940
rect 19628 23886 19630 23938
rect 19682 23886 20078 23938
rect 20130 23886 20132 23938
rect 19628 23884 20132 23886
rect 19628 23874 19684 23884
rect 20076 23874 20132 23884
rect 20188 23940 20244 23950
rect 20636 23940 20692 25566
rect 20188 23938 20692 23940
rect 20188 23886 20190 23938
rect 20242 23886 20692 23938
rect 20188 23884 20692 23886
rect 20748 24052 20804 24062
rect 20972 24052 21028 37996
rect 21420 37986 21476 37996
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 23212 28308 23268 28318
rect 21868 26964 21924 26974
rect 21308 26962 21924 26964
rect 21308 26910 21870 26962
rect 21922 26910 21924 26962
rect 21308 26908 21924 26910
rect 21084 26180 21140 26190
rect 21084 26178 21252 26180
rect 21084 26126 21086 26178
rect 21138 26126 21252 26178
rect 21084 26124 21252 26126
rect 21084 26114 21140 26124
rect 21196 25508 21252 26124
rect 21308 25730 21364 26908
rect 21868 26898 21924 26908
rect 22092 26964 22148 26974
rect 22092 26870 22148 26908
rect 22204 26962 22260 26974
rect 22204 26910 22206 26962
rect 22258 26910 22260 26962
rect 21308 25678 21310 25730
rect 21362 25678 21364 25730
rect 21308 25666 21364 25678
rect 21420 25730 21476 25742
rect 21420 25678 21422 25730
rect 21474 25678 21476 25730
rect 21420 25508 21476 25678
rect 21868 25508 21924 25518
rect 21196 25452 21476 25508
rect 21756 25506 21924 25508
rect 21756 25454 21870 25506
rect 21922 25454 21924 25506
rect 21756 25452 21924 25454
rect 21532 25394 21588 25406
rect 21532 25342 21534 25394
rect 21586 25342 21588 25394
rect 20972 23996 21476 24052
rect 20188 23874 20244 23884
rect 19964 23716 20020 23754
rect 19964 23650 20020 23660
rect 20412 23716 20468 23726
rect 20412 23714 20580 23716
rect 20412 23662 20414 23714
rect 20466 23662 20580 23714
rect 20412 23660 20580 23662
rect 20412 23650 20468 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23044 20244 23054
rect 20188 23042 20356 23044
rect 20188 22990 20190 23042
rect 20242 22990 20356 23042
rect 20188 22988 20356 22990
rect 20188 22978 20244 22988
rect 19628 22258 19684 22270
rect 19628 22206 19630 22258
rect 19682 22206 19684 22258
rect 19628 22148 19684 22206
rect 19740 22260 19796 22270
rect 19740 22166 19796 22204
rect 19964 22260 20020 22270
rect 19964 22166 20020 22204
rect 19628 21924 19684 22092
rect 20188 22148 20244 22158
rect 20188 22054 20244 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20300 21924 20356 22988
rect 19836 21914 20100 21924
rect 19628 21858 19684 21868
rect 20188 21868 20356 21924
rect 20412 22148 20468 22158
rect 20188 21812 20244 21868
rect 20412 21812 20468 22092
rect 19964 21756 20244 21812
rect 20300 21756 20468 21812
rect 20524 22146 20580 23660
rect 20524 22094 20526 22146
rect 20578 22094 20580 22146
rect 20524 21812 20580 22094
rect 19964 20914 20020 21756
rect 20300 21700 20356 21756
rect 20524 21746 20580 21756
rect 19964 20862 19966 20914
rect 20018 20862 20020 20914
rect 19964 20850 20020 20862
rect 20076 21644 20356 21700
rect 19628 20804 19684 20814
rect 19516 20802 19684 20804
rect 19516 20750 19630 20802
rect 19682 20750 19684 20802
rect 19516 20748 19684 20750
rect 19516 19908 19572 20748
rect 19628 20738 19684 20748
rect 20076 20802 20132 21644
rect 20748 21476 20804 23996
rect 21420 23044 21476 23996
rect 21532 23716 21588 25342
rect 21532 23650 21588 23660
rect 21420 22258 21476 22988
rect 21420 22206 21422 22258
rect 21474 22206 21476 22258
rect 21420 22194 21476 22206
rect 21532 22260 21588 22270
rect 21756 22260 21812 25452
rect 21868 25442 21924 25452
rect 22092 25506 22148 25518
rect 22092 25454 22094 25506
rect 22146 25454 22148 25506
rect 21532 22258 21812 22260
rect 21532 22206 21534 22258
rect 21586 22206 21812 22258
rect 21532 22204 21812 22206
rect 22092 23716 22148 25454
rect 22204 24948 22260 26910
rect 23212 26964 23268 28252
rect 24556 28308 24612 37998
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 24556 28242 24612 28252
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 22204 23940 22260 24892
rect 22428 26180 22484 26190
rect 22428 25508 22484 26124
rect 23212 26178 23268 26908
rect 25564 26404 25620 26414
rect 25564 26310 25620 26348
rect 37884 26404 37940 26414
rect 23212 26126 23214 26178
rect 23266 26126 23268 26178
rect 23212 26114 23268 26126
rect 25340 26290 25396 26302
rect 25340 26238 25342 26290
rect 25394 26238 25396 26290
rect 22764 25508 22820 25518
rect 22428 25506 22820 25508
rect 22428 25454 22766 25506
rect 22818 25454 22820 25506
rect 22428 25452 22820 25454
rect 22428 24724 22484 25452
rect 22764 25442 22820 25452
rect 23548 25396 23604 25406
rect 23548 25394 23828 25396
rect 23548 25342 23550 25394
rect 23602 25342 23828 25394
rect 23548 25340 23828 25342
rect 23548 25330 23604 25340
rect 23772 24946 23828 25340
rect 25340 25284 25396 26238
rect 37660 26290 37716 26302
rect 37660 26238 37662 26290
rect 37714 26238 37716 26290
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 25788 25284 25844 25294
rect 26236 25284 26292 25294
rect 25340 25282 26292 25284
rect 25340 25230 25790 25282
rect 25842 25230 26238 25282
rect 26290 25230 26292 25282
rect 25340 25228 26292 25230
rect 23772 24894 23774 24946
rect 23826 24894 23828 24946
rect 23772 24882 23828 24894
rect 25788 24836 25844 25228
rect 25788 24770 25844 24780
rect 22428 24052 22484 24668
rect 23324 24722 23380 24734
rect 23324 24670 23326 24722
rect 23378 24670 23380 24722
rect 23324 24052 23380 24670
rect 23996 24722 24052 24734
rect 23996 24670 23998 24722
rect 24050 24670 24052 24722
rect 23772 24612 23828 24622
rect 23660 24498 23716 24510
rect 23660 24446 23662 24498
rect 23714 24446 23716 24498
rect 22428 24050 22708 24052
rect 22428 23998 22430 24050
rect 22482 23998 22708 24050
rect 22428 23996 22708 23998
rect 23324 23996 23604 24052
rect 22428 23986 22484 23996
rect 22204 23874 22260 23884
rect 21196 22148 21252 22158
rect 21196 22054 21252 22092
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 20188 21420 20804 21476
rect 21532 21812 21588 22204
rect 19852 20692 19908 20702
rect 19852 20598 19908 20636
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20076 20244 20132 20254
rect 19740 20020 19796 20030
rect 19740 19926 19796 19964
rect 19516 19842 19572 19852
rect 20076 19684 20132 20188
rect 20188 20132 20244 21420
rect 21532 20916 21588 21756
rect 21532 20850 21588 20860
rect 21308 20804 21364 20814
rect 21308 20710 21364 20748
rect 20300 20690 20356 20702
rect 20300 20638 20302 20690
rect 20354 20638 20356 20690
rect 20300 20580 20356 20638
rect 21644 20580 21700 20590
rect 20300 20578 21812 20580
rect 20300 20526 21646 20578
rect 21698 20526 21812 20578
rect 20300 20524 21812 20526
rect 21644 20514 21700 20524
rect 20860 20132 20916 20142
rect 20188 19906 20244 20076
rect 20524 20076 20860 20132
rect 20188 19854 20190 19906
rect 20242 19854 20244 19906
rect 20188 19842 20244 19854
rect 20300 20018 20356 20030
rect 20300 19966 20302 20018
rect 20354 19966 20356 20018
rect 20076 19628 20244 19684
rect 19404 19404 19684 19460
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 18956 19012 19012 19182
rect 18956 18946 19012 18956
rect 19068 19346 19124 19358
rect 19068 19294 19070 19346
rect 19122 19294 19124 19346
rect 18956 18788 19012 18798
rect 19068 18788 19124 19294
rect 19404 19234 19460 19246
rect 19404 19182 19406 19234
rect 19458 19182 19460 19234
rect 19404 18900 19460 19182
rect 19404 18834 19460 18844
rect 19012 18732 19124 18788
rect 19180 18732 19348 18788
rect 18620 18622 18622 18674
rect 18674 18622 18676 18674
rect 18620 18610 18676 18622
rect 18732 18676 18788 18686
rect 18508 18498 18564 18508
rect 18732 18562 18788 18620
rect 18732 18510 18734 18562
rect 18786 18510 18788 18562
rect 18732 18498 18788 18510
rect 18956 18564 19012 18732
rect 19180 18676 19236 18732
rect 19180 18610 19236 18620
rect 19068 18564 19124 18574
rect 18956 18562 19124 18564
rect 18956 18510 19070 18562
rect 19122 18510 19124 18562
rect 18956 18508 19124 18510
rect 19068 18498 19124 18508
rect 18396 18450 18452 18462
rect 18396 18398 18398 18450
rect 18450 18398 18452 18450
rect 18396 18340 18452 18398
rect 18396 18274 18452 18284
rect 18956 18340 19012 18350
rect 18284 17838 18286 17890
rect 18338 17838 18340 17890
rect 18284 17826 18340 17838
rect 18844 18116 18900 18126
rect 18844 17890 18900 18060
rect 18844 17838 18846 17890
rect 18898 17838 18900 17890
rect 18844 17826 18900 17838
rect 18956 17892 19012 18284
rect 18956 17836 19124 17892
rect 17724 17378 17780 17388
rect 18396 17666 18452 17678
rect 18396 17614 18398 17666
rect 18450 17614 18452 17666
rect 18396 17108 18452 17614
rect 18956 17668 19012 17678
rect 18508 17108 18564 17118
rect 18396 17052 18508 17108
rect 18508 17042 18564 17052
rect 18956 15986 19012 17612
rect 19068 17666 19124 17836
rect 19068 17614 19070 17666
rect 19122 17614 19124 17666
rect 19068 17602 19124 17614
rect 19180 17554 19236 17566
rect 19180 17502 19182 17554
rect 19234 17502 19236 17554
rect 19068 17108 19124 17118
rect 19068 16098 19124 17052
rect 19180 16996 19236 17502
rect 19180 16930 19236 16940
rect 19068 16046 19070 16098
rect 19122 16046 19124 16098
rect 19068 16034 19124 16046
rect 18956 15934 18958 15986
rect 19010 15934 19012 15986
rect 18956 15922 19012 15934
rect 19292 15988 19348 18732
rect 19628 18676 19684 19404
rect 19964 19236 20020 19246
rect 19964 19010 20020 19180
rect 19964 18958 19966 19010
rect 20018 18958 20020 19010
rect 19964 18946 20020 18958
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18620 19796 18676
rect 19516 18564 19572 18574
rect 19516 18452 19572 18508
rect 19628 18452 19684 18462
rect 19516 18450 19684 18452
rect 19516 18398 19630 18450
rect 19682 18398 19684 18450
rect 19516 18396 19684 18398
rect 19628 18386 19684 18396
rect 19628 18228 19684 18238
rect 19628 17890 19684 18172
rect 19628 17838 19630 17890
rect 19682 17838 19684 17890
rect 19628 17826 19684 17838
rect 19404 17668 19460 17678
rect 19404 17574 19460 17612
rect 19740 17444 19796 18620
rect 20076 18450 20132 18462
rect 20076 18398 20078 18450
rect 20130 18398 20132 18450
rect 20076 18340 20132 18398
rect 20076 18274 20132 18284
rect 20188 17890 20244 19628
rect 20300 19348 20356 19966
rect 20300 19282 20356 19292
rect 20412 19124 20468 19134
rect 20412 19030 20468 19068
rect 20188 17838 20190 17890
rect 20242 17838 20244 17890
rect 20188 17826 20244 17838
rect 20300 19012 20356 19022
rect 20300 17892 20356 18956
rect 20524 17892 20580 20076
rect 20860 20038 20916 20076
rect 21196 19908 21252 19918
rect 21252 19852 21364 19908
rect 21196 19842 21252 19852
rect 20636 19348 20692 19358
rect 20636 18340 20692 19292
rect 20748 19010 20804 19022
rect 20748 18958 20750 19010
rect 20802 18958 20804 19010
rect 20748 18564 20804 18958
rect 20748 18470 20804 18508
rect 21196 18564 21252 18574
rect 20636 18274 20692 18284
rect 20300 17798 20356 17836
rect 20412 17836 20580 17892
rect 21084 18226 21140 18238
rect 21084 18174 21086 18226
rect 21138 18174 21140 18226
rect 20412 17668 20468 17836
rect 21084 17780 21140 18174
rect 21196 17892 21252 18508
rect 21308 18338 21364 19852
rect 21420 19906 21476 19918
rect 21420 19854 21422 19906
rect 21474 19854 21476 19906
rect 21420 19236 21476 19854
rect 21420 19234 21700 19236
rect 21420 19182 21422 19234
rect 21474 19182 21700 19234
rect 21420 19180 21700 19182
rect 21420 19170 21476 19180
rect 21420 18452 21476 18490
rect 21420 18386 21476 18396
rect 21308 18286 21310 18338
rect 21362 18286 21364 18338
rect 21308 18274 21364 18286
rect 21532 17892 21588 17902
rect 21196 17836 21476 17892
rect 20860 17724 21140 17780
rect 20524 17668 20580 17678
rect 20412 17666 20580 17668
rect 20412 17614 20526 17666
rect 20578 17614 20580 17666
rect 20412 17612 20580 17614
rect 20524 17602 20580 17612
rect 19628 17388 19796 17444
rect 20636 17556 20692 17566
rect 20860 17556 20916 17724
rect 20636 17554 20916 17556
rect 20636 17502 20638 17554
rect 20690 17502 20916 17554
rect 20636 17500 20916 17502
rect 21420 17554 21476 17836
rect 21532 17666 21588 17836
rect 21532 17614 21534 17666
rect 21586 17614 21588 17666
rect 21532 17602 21588 17614
rect 21420 17502 21422 17554
rect 21474 17502 21476 17554
rect 19292 15932 19572 15988
rect 18732 15876 18788 15886
rect 18508 15874 18788 15876
rect 18508 15822 18734 15874
rect 18786 15822 18788 15874
rect 18508 15820 18788 15822
rect 18060 15540 18116 15550
rect 17500 15538 18116 15540
rect 17500 15486 17502 15538
rect 17554 15486 18062 15538
rect 18114 15486 18116 15538
rect 17500 15484 18116 15486
rect 17500 15474 17556 15484
rect 18060 15474 18116 15484
rect 18284 15426 18340 15438
rect 18284 15374 18286 15426
rect 18338 15374 18340 15426
rect 17388 15202 17444 15214
rect 17388 15150 17390 15202
rect 17442 15150 17444 15202
rect 17388 15148 17444 15150
rect 16716 15092 17444 15148
rect 17724 15204 17780 15242
rect 17724 15138 17780 15148
rect 18172 15202 18228 15214
rect 18172 15150 18174 15202
rect 18226 15150 18228 15202
rect 16716 14642 16772 15092
rect 18172 14756 18228 15150
rect 16716 14590 16718 14642
rect 16770 14590 16772 14642
rect 16716 14578 16772 14590
rect 16828 14700 18228 14756
rect 15932 14438 15988 14476
rect 16828 13858 16884 14700
rect 16828 13806 16830 13858
rect 16882 13806 16884 13858
rect 16828 13794 16884 13806
rect 17388 14532 17444 14542
rect 17388 13748 17444 14476
rect 18172 14308 18228 14318
rect 18172 13858 18228 14252
rect 18172 13806 18174 13858
rect 18226 13806 18228 13858
rect 18172 13794 18228 13806
rect 17388 13654 17444 13692
rect 16716 13524 16772 13534
rect 15932 13522 16772 13524
rect 15932 13470 16718 13522
rect 16770 13470 16772 13522
rect 15932 13468 16772 13470
rect 15932 13074 15988 13468
rect 16716 13458 16772 13468
rect 15932 13022 15934 13074
rect 15986 13022 15988 13074
rect 15932 13010 15988 13022
rect 18060 13076 18116 13086
rect 18284 13076 18340 15374
rect 18508 15314 18564 15820
rect 18732 15810 18788 15820
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18508 14644 18564 15262
rect 18732 15428 18788 15438
rect 18732 15314 18788 15372
rect 19180 15428 19236 15438
rect 19180 15334 19236 15372
rect 18732 15262 18734 15314
rect 18786 15262 18788 15314
rect 18732 15250 18788 15262
rect 19404 15314 19460 15326
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 19292 15204 19348 15242
rect 19292 15138 19348 15148
rect 19404 14756 19460 15262
rect 19516 15316 19572 15932
rect 19628 15540 19684 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15484 19796 15540
rect 19628 15316 19684 15326
rect 19516 15314 19684 15316
rect 19516 15262 19630 15314
rect 19682 15262 19684 15314
rect 19516 15260 19684 15262
rect 19628 15250 19684 15260
rect 19740 15148 19796 15484
rect 20636 15316 20692 17500
rect 21420 17490 21476 17502
rect 21196 17442 21252 17454
rect 21196 17390 21198 17442
rect 21250 17390 21252 17442
rect 21196 17108 21252 17390
rect 21196 17042 21252 17052
rect 21532 17444 21588 17454
rect 21532 15428 21588 17388
rect 21644 16884 21700 19180
rect 21756 17780 21812 20524
rect 21980 20578 22036 20590
rect 21980 20526 21982 20578
rect 22034 20526 22036 20578
rect 21980 20356 22036 20526
rect 22092 20356 22148 23660
rect 22652 23380 22708 23996
rect 22764 23940 22820 23950
rect 22764 23846 22820 23884
rect 23100 23828 23156 23838
rect 23436 23828 23492 23838
rect 23100 23734 23156 23772
rect 23212 23826 23492 23828
rect 23212 23774 23438 23826
rect 23490 23774 23492 23826
rect 23212 23772 23492 23774
rect 22764 23380 22820 23390
rect 22652 23378 22820 23380
rect 22652 23326 22766 23378
rect 22818 23326 22820 23378
rect 22652 23324 22820 23326
rect 22764 23314 22820 23324
rect 22316 23044 22372 23054
rect 23212 23044 23268 23772
rect 23436 23762 23492 23772
rect 23548 23604 23604 23996
rect 23660 23714 23716 24446
rect 23772 23938 23828 24556
rect 23996 24052 24052 24670
rect 23996 23986 24052 23996
rect 24668 24724 24724 24734
rect 23772 23886 23774 23938
rect 23826 23886 23828 23938
rect 23772 23874 23828 23886
rect 23884 23938 23940 23950
rect 23884 23886 23886 23938
rect 23938 23886 23940 23938
rect 23660 23662 23662 23714
rect 23714 23662 23716 23714
rect 23660 23650 23716 23662
rect 22316 22950 22372 22988
rect 22764 22988 23268 23044
rect 23436 23548 23604 23604
rect 22764 22370 22820 22988
rect 22764 22318 22766 22370
rect 22818 22318 22820 22370
rect 22764 22306 22820 22318
rect 22204 22260 22260 22270
rect 22204 20802 22260 22204
rect 22204 20750 22206 20802
rect 22258 20750 22260 20802
rect 22204 20738 22260 20750
rect 22428 22258 22484 22270
rect 22428 22206 22430 22258
rect 22482 22206 22484 22258
rect 22428 20580 22484 22206
rect 22540 22260 22596 22270
rect 22540 22166 22596 22204
rect 23212 22148 23268 22158
rect 23212 20914 23268 22092
rect 23212 20862 23214 20914
rect 23266 20862 23268 20914
rect 23212 20850 23268 20862
rect 23436 21474 23492 23548
rect 23884 22148 23940 23886
rect 23884 22082 23940 22092
rect 24332 23940 24388 23950
rect 24332 21812 24388 23884
rect 24668 23604 24724 24668
rect 25228 24724 25284 24734
rect 25228 24630 25284 24668
rect 26012 24612 26068 24622
rect 25340 24610 26068 24612
rect 25340 24558 26014 24610
rect 26066 24558 26068 24610
rect 25340 24556 26068 24558
rect 25228 24052 25284 24062
rect 25340 24052 25396 24556
rect 26012 24546 26068 24556
rect 25228 24050 25396 24052
rect 25228 23998 25230 24050
rect 25282 23998 25396 24050
rect 25228 23996 25396 23998
rect 25228 23986 25284 23996
rect 25116 23940 25172 23978
rect 25116 23874 25172 23884
rect 25788 23940 25844 23950
rect 26124 23940 26180 23950
rect 25788 23938 26180 23940
rect 25788 23886 25790 23938
rect 25842 23886 26126 23938
rect 26178 23886 26180 23938
rect 25788 23884 26180 23886
rect 25788 23874 25844 23884
rect 26124 23874 26180 23884
rect 26236 23940 26292 25228
rect 26572 25284 26628 25294
rect 26572 25190 26628 25228
rect 37660 25284 37716 26238
rect 37884 25506 37940 26348
rect 39900 26178 39956 26190
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 25620 39956 26126
rect 39900 25554 39956 25564
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37884 25454 37886 25506
rect 37938 25454 37940 25506
rect 37884 25442 37940 25454
rect 37660 25218 37716 25228
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 37660 24724 37716 24734
rect 37660 24630 37716 24668
rect 26236 23874 26292 23884
rect 26348 24612 26404 24622
rect 25564 23828 25620 23838
rect 25452 23772 25564 23828
rect 25340 23716 25396 23726
rect 25340 23622 25396 23660
rect 24668 23538 24724 23548
rect 25228 23548 25284 23558
rect 25228 22596 25284 23492
rect 25004 22540 25284 22596
rect 24892 22484 24948 22494
rect 25004 22484 25060 22540
rect 24892 22482 25060 22484
rect 24892 22430 24894 22482
rect 24946 22430 25060 22482
rect 24892 22428 25060 22430
rect 24892 22418 24948 22428
rect 23436 21422 23438 21474
rect 23490 21422 23492 21474
rect 22428 20514 22484 20524
rect 23100 20690 23156 20702
rect 23100 20638 23102 20690
rect 23154 20638 23156 20690
rect 23100 20580 23156 20638
rect 23100 20514 23156 20524
rect 23324 20578 23380 20590
rect 23324 20526 23326 20578
rect 23378 20526 23380 20578
rect 22092 20300 22596 20356
rect 21980 18676 22036 20300
rect 22092 20132 22148 20142
rect 22092 19348 22148 20076
rect 22092 19346 22372 19348
rect 22092 19294 22094 19346
rect 22146 19294 22372 19346
rect 22092 19292 22372 19294
rect 22092 19282 22148 19292
rect 21980 18610 22036 18620
rect 22316 18674 22372 19292
rect 22316 18622 22318 18674
rect 22370 18622 22372 18674
rect 22316 18610 22372 18622
rect 21868 18564 21924 18574
rect 21868 18470 21924 18508
rect 22428 18564 22484 18574
rect 22428 18470 22484 18508
rect 21980 18450 22036 18462
rect 21980 18398 21982 18450
rect 22034 18398 22036 18450
rect 21868 18228 21924 18238
rect 21868 18134 21924 18172
rect 21756 17714 21812 17724
rect 21868 17892 21924 17902
rect 21868 17778 21924 17836
rect 21980 17892 22036 18398
rect 22540 18228 22596 20300
rect 23324 18676 23380 20526
rect 23436 20132 23492 21422
rect 23772 21810 24388 21812
rect 23772 21758 24334 21810
rect 24386 21758 24388 21810
rect 23772 21756 24388 21758
rect 23772 20802 23828 21756
rect 24332 21746 24388 21756
rect 23772 20750 23774 20802
rect 23826 20750 23828 20802
rect 23436 20076 23716 20132
rect 23548 18676 23604 18686
rect 22540 18162 22596 18172
rect 22876 18674 23604 18676
rect 22876 18622 23550 18674
rect 23602 18622 23604 18674
rect 22876 18620 23604 18622
rect 22652 17892 22708 17902
rect 21980 17890 22708 17892
rect 21980 17838 21982 17890
rect 22034 17838 22654 17890
rect 22706 17838 22708 17890
rect 21980 17836 22708 17838
rect 21980 17826 22036 17836
rect 22652 17826 22708 17836
rect 21868 17726 21870 17778
rect 21922 17726 21924 17778
rect 21868 17714 21924 17726
rect 22876 17554 22932 18620
rect 23436 18452 23492 18620
rect 23548 18610 23604 18620
rect 23660 18452 23716 20076
rect 23772 19684 23828 20750
rect 24108 21586 24164 21598
rect 24108 21534 24110 21586
rect 24162 21534 24164 21586
rect 23996 20690 24052 20702
rect 23996 20638 23998 20690
rect 24050 20638 24052 20690
rect 23996 20356 24052 20638
rect 24108 20580 24164 21534
rect 25228 21586 25284 22540
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 25228 21522 25284 21534
rect 24556 21476 24612 21486
rect 24220 21028 24276 21038
rect 24220 20934 24276 20972
rect 24444 20916 24500 20926
rect 24444 20822 24500 20860
rect 24556 20914 24612 21420
rect 24556 20862 24558 20914
rect 24610 20862 24612 20914
rect 24556 20850 24612 20862
rect 24668 20692 24724 20702
rect 24668 20598 24724 20636
rect 24108 20514 24164 20524
rect 23996 20290 24052 20300
rect 25452 20244 25508 23772
rect 25564 23762 25620 23772
rect 26348 23826 26404 24556
rect 28140 24612 28196 24622
rect 28140 24518 28196 24556
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23940 37716 23950
rect 37660 23846 37716 23884
rect 26348 23774 26350 23826
rect 26402 23774 26404 23826
rect 26348 23762 26404 23774
rect 26460 23828 26516 23838
rect 26460 23734 26516 23772
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37660 22370 37716 22382
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 37660 21812 37716 22318
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 37660 21746 37716 21756
rect 28812 21700 28868 21710
rect 28812 21606 28868 21644
rect 28588 21588 28644 21598
rect 28140 21532 28588 21588
rect 26012 21476 26068 21486
rect 26012 21382 26068 21420
rect 27020 21476 27076 21486
rect 27020 20914 27076 21420
rect 28140 21476 28196 21532
rect 28588 21494 28644 21532
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21588 40068 21598
rect 28140 21382 28196 21420
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 27020 20862 27022 20914
rect 27074 20862 27076 20914
rect 27020 20850 27076 20862
rect 40012 20914 40068 20926
rect 40012 20862 40014 20914
rect 40066 20862 40068 20914
rect 37660 20802 37716 20814
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 26012 20690 26068 20702
rect 26012 20638 26014 20690
rect 26066 20638 26068 20690
rect 26012 20580 26068 20638
rect 26908 20692 26964 20702
rect 26908 20598 26964 20636
rect 25452 20178 25508 20188
rect 25788 20524 26068 20580
rect 26124 20580 26180 20590
rect 26124 20578 26292 20580
rect 26124 20526 26126 20578
rect 26178 20526 26292 20578
rect 26124 20524 26292 20526
rect 25788 20132 25844 20524
rect 26124 20514 26180 20524
rect 25564 20076 25844 20132
rect 25900 20356 25956 20366
rect 25452 20018 25508 20030
rect 25452 19966 25454 20018
rect 25506 19966 25508 20018
rect 23772 19618 23828 19628
rect 24780 19908 24836 19918
rect 25452 19908 25508 19966
rect 24780 19906 25508 19908
rect 24780 19854 24782 19906
rect 24834 19854 25508 19906
rect 24780 19852 25508 19854
rect 24220 19346 24276 19358
rect 24220 19294 24222 19346
rect 24274 19294 24276 19346
rect 23436 18386 23492 18396
rect 23548 18396 23716 18452
rect 23772 19124 23828 19134
rect 23772 18450 23828 19068
rect 24220 19124 24276 19294
rect 24220 19058 24276 19068
rect 23772 18398 23774 18450
rect 23826 18398 23828 18450
rect 22988 17780 23044 17790
rect 22988 17778 23492 17780
rect 22988 17726 22990 17778
rect 23042 17726 23492 17778
rect 22988 17724 23492 17726
rect 22988 17714 23044 17724
rect 22876 17502 22878 17554
rect 22930 17502 22932 17554
rect 22876 17490 22932 17502
rect 21756 16884 21812 16894
rect 21644 16828 21756 16884
rect 21756 16770 21812 16828
rect 21756 16718 21758 16770
rect 21810 16718 21812 16770
rect 21756 15540 21812 16718
rect 23212 16100 23268 16110
rect 23212 16006 23268 16044
rect 23436 16098 23492 17724
rect 23548 16882 23604 18396
rect 23772 18386 23828 18398
rect 24780 17444 24836 19852
rect 25228 19684 25284 19694
rect 25116 19236 25172 19246
rect 25116 19142 25172 19180
rect 25228 18450 25284 19628
rect 25452 19348 25508 19358
rect 25564 19348 25620 20076
rect 25452 19346 25620 19348
rect 25452 19294 25454 19346
rect 25506 19294 25620 19346
rect 25452 19292 25620 19294
rect 25788 19908 25844 19918
rect 25452 19282 25508 19292
rect 25788 19234 25844 19852
rect 25788 19182 25790 19234
rect 25842 19182 25844 19234
rect 25788 19170 25844 19182
rect 25564 19124 25620 19134
rect 25564 19030 25620 19068
rect 25228 18398 25230 18450
rect 25282 18398 25284 18450
rect 25228 17780 25284 18398
rect 25340 19010 25396 19022
rect 25340 18958 25342 19010
rect 25394 18958 25396 19010
rect 25340 18452 25396 18958
rect 25900 18674 25956 20300
rect 26236 20130 26292 20524
rect 26236 20078 26238 20130
rect 26290 20078 26292 20130
rect 26236 20066 26292 20078
rect 28364 19908 28420 19918
rect 28364 19814 28420 19852
rect 37660 19908 37716 20750
rect 40012 20244 40068 20862
rect 40012 20178 40068 20188
rect 37660 19842 37716 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 25900 18622 25902 18674
rect 25954 18622 25956 18674
rect 25900 18610 25956 18622
rect 26348 19124 26404 19134
rect 25340 18386 25396 18396
rect 25676 18452 25732 18462
rect 25676 18358 25732 18396
rect 26124 18452 26180 18462
rect 26124 18358 26180 18396
rect 25452 18340 25508 18350
rect 25452 18246 25508 18284
rect 26012 18338 26068 18350
rect 26012 18286 26014 18338
rect 26066 18286 26068 18338
rect 25900 17780 25956 17790
rect 26012 17780 26068 18286
rect 25228 17724 25508 17780
rect 25116 17666 25172 17678
rect 25116 17614 25118 17666
rect 25170 17614 25172 17666
rect 25116 17444 25172 17614
rect 24668 17442 25172 17444
rect 24668 17390 24782 17442
rect 24834 17390 25172 17442
rect 24668 17388 25172 17390
rect 23548 16830 23550 16882
rect 23602 16830 23604 16882
rect 23548 16818 23604 16830
rect 24332 16884 24388 16894
rect 24332 16212 24388 16828
rect 24668 16212 24724 17388
rect 24780 17378 24836 17388
rect 25228 17108 25284 17118
rect 25228 17014 25284 17052
rect 25452 17106 25508 17724
rect 25900 17778 26068 17780
rect 25900 17726 25902 17778
rect 25954 17726 26068 17778
rect 25900 17724 26068 17726
rect 25900 17714 25956 17724
rect 25452 17054 25454 17106
rect 25506 17054 25508 17106
rect 25452 17042 25508 17054
rect 26012 16994 26068 17006
rect 26012 16942 26014 16994
rect 26066 16942 26068 16994
rect 25900 16884 25956 16894
rect 26012 16884 26068 16942
rect 26236 16996 26292 17006
rect 26236 16902 26292 16940
rect 26348 16994 26404 19068
rect 27020 18452 27076 18462
rect 27020 17106 27076 18396
rect 37660 18450 37716 18462
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 28028 17778 28084 17790
rect 28028 17726 28030 17778
rect 28082 17726 28084 17778
rect 27020 17054 27022 17106
rect 27074 17054 27076 17106
rect 27020 17042 27076 17054
rect 27132 17108 27188 17118
rect 26348 16942 26350 16994
rect 26402 16942 26404 16994
rect 25900 16882 26068 16884
rect 25900 16830 25902 16882
rect 25954 16830 26068 16882
rect 25900 16828 26068 16830
rect 25900 16818 25956 16828
rect 24332 16210 24724 16212
rect 24332 16158 24334 16210
rect 24386 16158 24724 16210
rect 24332 16156 24724 16158
rect 25340 16770 25396 16782
rect 25340 16718 25342 16770
rect 25394 16718 25396 16770
rect 25340 16212 25396 16718
rect 25452 16212 25508 16222
rect 25340 16210 25508 16212
rect 25340 16158 25454 16210
rect 25506 16158 25508 16210
rect 25340 16156 25508 16158
rect 24332 16146 24388 16156
rect 23436 16046 23438 16098
rect 23490 16046 23492 16098
rect 21756 15484 22036 15540
rect 20972 15316 21028 15326
rect 20636 15314 21028 15316
rect 20636 15262 20974 15314
rect 21026 15262 21028 15314
rect 20636 15260 21028 15262
rect 20972 15250 21028 15260
rect 21196 15316 21252 15326
rect 21196 15222 21252 15260
rect 21532 15314 21588 15372
rect 21532 15262 21534 15314
rect 21586 15262 21588 15314
rect 21532 15250 21588 15262
rect 21644 15314 21700 15326
rect 21644 15262 21646 15314
rect 21698 15262 21700 15314
rect 19516 15092 19796 15148
rect 19964 15204 20020 15214
rect 19516 14868 19572 15092
rect 19516 14812 19684 14868
rect 19180 14700 19460 14756
rect 18732 14644 18788 14654
rect 18508 14588 18732 14644
rect 18732 14578 18788 14588
rect 18844 14644 18900 14654
rect 19180 14644 19236 14700
rect 18844 14642 19236 14644
rect 18844 14590 18846 14642
rect 18898 14590 19236 14642
rect 18844 14588 19236 14590
rect 19516 14644 19572 14654
rect 18060 13074 18340 13076
rect 18060 13022 18062 13074
rect 18114 13022 18340 13074
rect 18060 13020 18340 13022
rect 18620 13748 18676 13758
rect 18620 13186 18676 13692
rect 18620 13134 18622 13186
rect 18674 13134 18676 13186
rect 18620 13074 18676 13134
rect 18620 13022 18622 13074
rect 18674 13022 18676 13074
rect 15148 12910 15150 12962
rect 15202 12910 15204 12962
rect 15148 12898 15204 12910
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 18060 8428 18116 13020
rect 18620 13010 18676 13022
rect 17612 8372 18116 8428
rect 18844 8428 18900 14588
rect 19516 14550 19572 14588
rect 19292 14530 19348 14542
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 19292 14420 19348 14478
rect 19628 14420 19684 14812
rect 19964 14530 20020 15148
rect 21644 15204 21700 15262
rect 21868 15314 21924 15326
rect 21868 15262 21870 15314
rect 21922 15262 21924 15314
rect 21644 15138 21700 15148
rect 21756 15202 21812 15214
rect 21756 15150 21758 15202
rect 21810 15150 21812 15202
rect 20524 14644 20580 14654
rect 20748 14644 20804 14654
rect 20524 14642 20748 14644
rect 20524 14590 20526 14642
rect 20578 14590 20748 14642
rect 20524 14588 20748 14590
rect 20524 14578 20580 14588
rect 19964 14478 19966 14530
rect 20018 14478 20020 14530
rect 19964 14466 20020 14478
rect 19292 14364 19684 14420
rect 19740 14308 19796 14318
rect 19628 14306 19796 14308
rect 19628 14254 19742 14306
rect 19794 14254 19796 14306
rect 19628 14252 19796 14254
rect 19180 13186 19236 13198
rect 19180 13134 19182 13186
rect 19234 13134 19236 13186
rect 19180 13074 19236 13134
rect 19628 13188 19684 14252
rect 19740 14242 19796 14252
rect 19852 14308 19908 14346
rect 19852 14242 19908 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20748 13748 20804 14588
rect 21756 14420 21812 15150
rect 21420 14364 21812 14420
rect 21868 14420 21924 15262
rect 21980 14644 22036 15484
rect 23436 15316 23492 16046
rect 23884 16100 23940 16110
rect 23884 16006 23940 16044
rect 24668 16098 24724 16156
rect 25452 16146 25508 16156
rect 24668 16046 24670 16098
rect 24722 16046 24724 16098
rect 24668 16034 24724 16046
rect 26348 16100 26404 16942
rect 27132 16994 27188 17052
rect 28028 17108 28084 17726
rect 28028 17042 28084 17052
rect 37660 17108 37716 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37660 17042 37716 17052
rect 27132 16942 27134 16994
rect 27186 16942 27188 16994
rect 27132 16930 27188 16942
rect 27580 16884 27636 16894
rect 27580 16210 27636 16828
rect 37660 16884 37716 16894
rect 37660 16790 37716 16828
rect 40012 16658 40068 16670
rect 40012 16606 40014 16658
rect 40066 16606 40068 16658
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 27580 16158 27582 16210
rect 27634 16158 27636 16210
rect 27580 16146 27636 16158
rect 40012 16212 40068 16606
rect 40012 16146 40068 16156
rect 26348 16034 26404 16044
rect 23548 15874 23604 15886
rect 23548 15822 23550 15874
rect 23602 15822 23604 15874
rect 23548 15540 23604 15822
rect 23660 15876 23716 15886
rect 23660 15782 23716 15820
rect 25788 15876 25844 15886
rect 23548 15484 23940 15540
rect 23884 15426 23940 15484
rect 23884 15374 23886 15426
rect 23938 15374 23940 15426
rect 23884 15362 23940 15374
rect 23436 15250 23492 15260
rect 23772 15092 23828 15102
rect 23660 15090 23828 15092
rect 23660 15038 23774 15090
rect 23826 15038 23828 15090
rect 23660 15036 23828 15038
rect 22092 14644 22148 14654
rect 21980 14588 22092 14644
rect 22092 14550 22148 14588
rect 22876 14644 22932 14654
rect 22876 14530 22932 14588
rect 23660 14642 23716 15036
rect 23772 15026 23828 15036
rect 23660 14590 23662 14642
rect 23714 14590 23716 14642
rect 23660 14578 23716 14590
rect 23996 14644 24052 14654
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 22876 14466 22932 14478
rect 22428 14420 22484 14430
rect 21868 14418 22484 14420
rect 21868 14366 22430 14418
rect 22482 14366 22484 14418
rect 21868 14364 22484 14366
rect 21420 13858 21476 14364
rect 22428 14354 22484 14364
rect 22540 14418 22596 14430
rect 22540 14366 22542 14418
rect 22594 14366 22596 14418
rect 21420 13806 21422 13858
rect 21474 13806 21476 13858
rect 21420 13794 21476 13806
rect 20748 13654 20804 13692
rect 19628 13122 19684 13132
rect 20300 13634 20356 13646
rect 20300 13582 20302 13634
rect 20354 13582 20356 13634
rect 19180 13022 19182 13074
rect 19234 13022 19236 13074
rect 19180 13010 19236 13022
rect 20300 12852 20356 13582
rect 22540 13524 22596 14366
rect 23996 13970 24052 14588
rect 23996 13918 23998 13970
rect 24050 13918 24052 13970
rect 23996 13906 24052 13918
rect 25788 14642 25844 15820
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 25788 14590 25790 14642
rect 25842 14590 25844 14642
rect 22540 13458 22596 13468
rect 23548 13634 23604 13646
rect 23548 13582 23550 13634
rect 23602 13582 23604 13634
rect 23548 13524 23604 13582
rect 23548 13458 23604 13468
rect 24556 13524 24612 13534
rect 20636 13188 20692 13198
rect 20636 13094 20692 13132
rect 20748 12852 20804 12862
rect 20300 12850 20804 12852
rect 20300 12798 20750 12850
rect 20802 12798 20804 12850
rect 20300 12796 20804 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20748 8428 20804 12796
rect 18844 8372 19124 8428
rect 20748 8372 21140 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17612 3554 17668 8372
rect 19068 4338 19124 8372
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4274 19124 4286
rect 18844 4116 18900 4126
rect 18620 3668 18676 3678
rect 17612 3502 17614 3554
rect 17666 3502 17668 3554
rect 17612 3490 17668 3502
rect 18172 3666 18676 3668
rect 18172 3614 18622 3666
rect 18674 3614 18676 3666
rect 18172 3612 18676 3614
rect 18172 800 18228 3612
rect 18620 3602 18676 3612
rect 18844 800 18900 4060
rect 20076 4116 20132 4126
rect 20076 4022 20132 4060
rect 20860 3668 20916 3678
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 3612
rect 21084 3554 21140 8372
rect 24220 4116 24276 4126
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 22876 3668 22932 3678
rect 21084 3502 21086 3554
rect 21138 3502 21140 3554
rect 21084 3490 21140 3502
rect 22876 800 22932 3612
rect 24220 800 24276 4060
rect 24556 3554 24612 13468
rect 25788 8428 25844 14590
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 25228 8372 25844 8428
rect 25228 4338 25284 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 20832 0 20944 800
rect 22848 0 22960 800
rect 24192 0 24304 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 14924 37996 14980 38052
rect 1708 36988 1764 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 13468 28476 13524 28532
rect 14588 28588 14644 28644
rect 4172 28252 4228 28308
rect 1932 27186 1988 27188
rect 1932 27134 1934 27186
rect 1934 27134 1986 27186
rect 1986 27134 1988 27186
rect 1932 27132 1988 27134
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 11228 27020 11284 27076
rect 13132 26908 13188 26964
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 13916 27132 13972 27188
rect 13804 27020 13860 27076
rect 13356 25676 13412 25732
rect 15932 38050 15988 38052
rect 15932 37998 15934 38050
rect 15934 37998 15986 38050
rect 15986 37998 15988 38050
rect 15932 37996 15988 37998
rect 16156 37436 16212 37492
rect 15484 36652 15540 36708
rect 16716 36706 16772 36708
rect 16716 36654 16718 36706
rect 16718 36654 16770 36706
rect 16770 36654 16772 36706
rect 16716 36652 16772 36654
rect 14924 28476 14980 28532
rect 14364 27468 14420 27524
rect 14252 26962 14308 26964
rect 14252 26910 14254 26962
rect 14254 26910 14306 26962
rect 14306 26910 14308 26962
rect 14252 26908 14308 26910
rect 14140 26124 14196 26180
rect 13916 25730 13972 25732
rect 13916 25678 13918 25730
rect 13918 25678 13970 25730
rect 13970 25678 13972 25730
rect 13916 25676 13972 25678
rect 12460 25228 12516 25284
rect 13468 24946 13524 24948
rect 13468 24894 13470 24946
rect 13470 24894 13522 24946
rect 13522 24894 13524 24946
rect 13468 24892 13524 24894
rect 16268 28642 16324 28644
rect 16268 28590 16270 28642
rect 16270 28590 16322 28642
rect 16322 28590 16324 28642
rect 16268 28588 16324 28590
rect 16828 28642 16884 28644
rect 16828 28590 16830 28642
rect 16830 28590 16882 28642
rect 16882 28590 16884 28642
rect 16828 28588 16884 28590
rect 15708 27468 15764 27524
rect 14924 27020 14980 27076
rect 15148 27132 15204 27188
rect 15596 27020 15652 27076
rect 15036 26962 15092 26964
rect 15036 26910 15038 26962
rect 15038 26910 15090 26962
rect 15090 26910 15092 26962
rect 15036 26908 15092 26910
rect 14476 26850 14532 26852
rect 14476 26798 14478 26850
rect 14478 26798 14530 26850
rect 14530 26798 14532 26850
rect 14476 26796 14532 26798
rect 15820 27020 15876 27076
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 22876 38220 22932 38276
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 20188 37436 20244 37492
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 17388 28476 17444 28532
rect 17276 26908 17332 26964
rect 18620 28530 18676 28532
rect 18620 28478 18622 28530
rect 18622 28478 18674 28530
rect 18674 28478 18676 28530
rect 18620 28476 18676 28478
rect 17948 27020 18004 27076
rect 15372 26796 15428 26852
rect 14028 25004 14084 25060
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 13692 23660 13748 23716
rect 13804 23938 13860 23940
rect 13804 23886 13806 23938
rect 13806 23886 13858 23938
rect 13858 23886 13860 23938
rect 13804 23884 13860 23886
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 22092 4228 22148
rect 11676 23042 11732 23044
rect 11676 22990 11678 23042
rect 11678 22990 11730 23042
rect 11730 22990 11732 23042
rect 11676 22988 11732 22990
rect 11004 21980 11060 22036
rect 13132 21980 13188 22036
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 9996 21532 10052 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1932 20860 1988 20916
rect 9996 20914 10052 20916
rect 9996 20862 9998 20914
rect 9998 20862 10050 20914
rect 10050 20862 10052 20914
rect 9996 20860 10052 20862
rect 13916 22876 13972 22932
rect 14364 23772 14420 23828
rect 14140 23660 14196 23716
rect 14252 23042 14308 23044
rect 14252 22990 14254 23042
rect 14254 22990 14306 23042
rect 14306 22990 14308 23042
rect 14252 22988 14308 22990
rect 14028 21980 14084 22036
rect 13916 21868 13972 21924
rect 14028 21644 14084 21700
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 15708 26178 15764 26180
rect 15708 26126 15710 26178
rect 15710 26126 15762 26178
rect 15762 26126 15764 26178
rect 15708 26124 15764 26126
rect 17724 26124 17780 26180
rect 15148 24892 15204 24948
rect 14588 23884 14644 23940
rect 15036 23772 15092 23828
rect 14924 22876 14980 22932
rect 15148 23660 15204 23716
rect 17500 24780 17556 24836
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19516 26178 19572 26180
rect 19516 26126 19518 26178
rect 19518 26126 19570 26178
rect 19570 26126 19572 26178
rect 19516 26124 19572 26126
rect 19964 26178 20020 26180
rect 19964 26126 19966 26178
rect 19966 26126 20018 26178
rect 20018 26126 20020 26178
rect 19964 26124 20020 26126
rect 20412 26124 20468 26180
rect 18172 24892 18228 24948
rect 15148 23266 15204 23268
rect 15148 23214 15150 23266
rect 15150 23214 15202 23266
rect 15202 23214 15204 23266
rect 15148 23212 15204 23214
rect 14588 22258 14644 22260
rect 14588 22206 14590 22258
rect 14590 22206 14642 22258
rect 14642 22206 14644 22258
rect 14588 22204 14644 22206
rect 14476 21980 14532 22036
rect 14476 21644 14532 21700
rect 13580 20802 13636 20804
rect 13580 20750 13582 20802
rect 13582 20750 13634 20802
rect 13634 20750 13636 20802
rect 13580 20748 13636 20750
rect 12124 20690 12180 20692
rect 12124 20638 12126 20690
rect 12126 20638 12178 20690
rect 12178 20638 12180 20690
rect 12124 20636 12180 20638
rect 12236 20524 12292 20580
rect 13804 20578 13860 20580
rect 13804 20526 13806 20578
rect 13806 20526 13858 20578
rect 13858 20526 13860 20578
rect 13804 20524 13860 20526
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 11452 18396 11508 18452
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 12012 17612 12068 17668
rect 1932 16828 1988 16884
rect 4284 16940 4340 16996
rect 11788 16940 11844 16996
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1932 16156 1988 16212
rect 14924 21698 14980 21700
rect 14924 21646 14926 21698
rect 14926 21646 14978 21698
rect 14978 21646 14980 21698
rect 14924 21644 14980 21646
rect 14700 20860 14756 20916
rect 15820 23212 15876 23268
rect 14812 20412 14868 20468
rect 14252 19180 14308 19236
rect 14364 19404 14420 19460
rect 14924 19404 14980 19460
rect 14924 19234 14980 19236
rect 14924 19182 14926 19234
rect 14926 19182 14978 19234
rect 14978 19182 14980 19234
rect 14924 19180 14980 19182
rect 18284 24834 18340 24836
rect 18284 24782 18286 24834
rect 18286 24782 18338 24834
rect 18338 24782 18340 24834
rect 18284 24780 18340 24782
rect 19292 24780 19348 24836
rect 17500 23714 17556 23716
rect 17500 23662 17502 23714
rect 17502 23662 17554 23714
rect 17554 23662 17556 23714
rect 17500 23660 17556 23662
rect 17836 23826 17892 23828
rect 17836 23774 17838 23826
rect 17838 23774 17890 23826
rect 17890 23774 17892 23826
rect 17836 23772 17892 23774
rect 17500 23042 17556 23044
rect 17500 22990 17502 23042
rect 17502 22990 17554 23042
rect 17554 22990 17556 23042
rect 17500 22988 17556 22990
rect 19404 23826 19460 23828
rect 19404 23774 19406 23826
rect 19406 23774 19458 23826
rect 19458 23774 19460 23826
rect 19404 23772 19460 23774
rect 16156 22370 16212 22372
rect 16156 22318 16158 22370
rect 16158 22318 16210 22370
rect 16210 22318 16212 22370
rect 16156 22316 16212 22318
rect 17612 22316 17668 22372
rect 15932 22258 15988 22260
rect 15932 22206 15934 22258
rect 15934 22206 15986 22258
rect 15986 22206 15988 22258
rect 15932 22204 15988 22206
rect 17164 22204 17220 22260
rect 15820 21868 15876 21924
rect 17388 22258 17444 22260
rect 17388 22206 17390 22258
rect 17390 22206 17442 22258
rect 17442 22206 17444 22258
rect 17388 22204 17444 22206
rect 18172 22988 18228 23044
rect 17164 21980 17220 22036
rect 16380 20860 16436 20916
rect 15708 20748 15764 20804
rect 15372 20690 15428 20692
rect 15372 20638 15374 20690
rect 15374 20638 15426 20690
rect 15426 20638 15428 20690
rect 15372 20636 15428 20638
rect 15260 20076 15316 20132
rect 16156 20802 16212 20804
rect 16156 20750 16158 20802
rect 16158 20750 16210 20802
rect 16210 20750 16212 20802
rect 16156 20748 16212 20750
rect 15484 19404 15540 19460
rect 17500 21980 17556 22036
rect 17724 21474 17780 21476
rect 17724 21422 17726 21474
rect 17726 21422 17778 21474
rect 17778 21422 17780 21474
rect 17724 21420 17780 21422
rect 17500 21308 17556 21364
rect 17164 20914 17220 20916
rect 17164 20862 17166 20914
rect 17166 20862 17218 20914
rect 17218 20862 17220 20914
rect 17164 20860 17220 20862
rect 17948 21026 18004 21028
rect 17948 20974 17950 21026
rect 17950 20974 18002 21026
rect 18002 20974 18004 21026
rect 17948 20972 18004 20974
rect 17388 20802 17444 20804
rect 17388 20750 17390 20802
rect 17390 20750 17442 20802
rect 17442 20750 17444 20802
rect 17388 20748 17444 20750
rect 18172 21308 18228 21364
rect 18508 22204 18564 22260
rect 18620 22092 18676 22148
rect 19292 21980 19348 22036
rect 18508 20748 18564 20804
rect 17724 20188 17780 20244
rect 18060 20130 18116 20132
rect 18060 20078 18062 20130
rect 18062 20078 18114 20130
rect 18114 20078 18116 20130
rect 18060 20076 18116 20078
rect 18620 21308 18676 21364
rect 18732 20636 18788 20692
rect 16156 19234 16212 19236
rect 16156 19182 16158 19234
rect 16158 19182 16210 19234
rect 16210 19182 16212 19234
rect 16156 19180 16212 19182
rect 17836 19346 17892 19348
rect 17836 19294 17838 19346
rect 17838 19294 17890 19346
rect 17890 19294 17892 19346
rect 17836 19292 17892 19294
rect 17052 19234 17108 19236
rect 17052 19182 17054 19234
rect 17054 19182 17106 19234
rect 17106 19182 17108 19234
rect 17052 19180 17108 19182
rect 18060 19234 18116 19236
rect 18060 19182 18062 19234
rect 18062 19182 18114 19234
rect 18114 19182 18116 19234
rect 18060 19180 18116 19182
rect 16380 19068 16436 19124
rect 17388 18844 17444 18900
rect 18060 18956 18116 19012
rect 16828 18732 16884 18788
rect 15036 18396 15092 18452
rect 14924 18284 14980 18340
rect 14924 17388 14980 17444
rect 14812 16940 14868 16996
rect 14476 16828 14532 16884
rect 14252 16098 14308 16100
rect 14252 16046 14254 16098
rect 14254 16046 14306 16098
rect 14306 16046 14308 16098
rect 14252 16044 14308 16046
rect 16492 18284 16548 18340
rect 17052 18284 17108 18340
rect 15484 17836 15540 17892
rect 15260 17666 15316 17668
rect 15260 17614 15262 17666
rect 15262 17614 15314 17666
rect 15314 17614 15316 17666
rect 15260 17612 15316 17614
rect 17724 18284 17780 18340
rect 17388 17612 17444 17668
rect 15484 17388 15540 17444
rect 15372 17106 15428 17108
rect 15372 17054 15374 17106
rect 15374 17054 15426 17106
rect 15426 17054 15428 17106
rect 15372 17052 15428 17054
rect 15148 16716 15204 16772
rect 15372 16828 15428 16884
rect 15932 16770 15988 16772
rect 15932 16718 15934 16770
rect 15934 16718 15986 16770
rect 15986 16718 15988 16770
rect 15932 16716 15988 16718
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 17948 18396 18004 18452
rect 17948 17890 18004 17892
rect 17948 17838 17950 17890
rect 17950 17838 18002 17890
rect 18002 17838 18004 17890
rect 17948 17836 18004 17838
rect 18284 18732 18340 18788
rect 19180 20412 19236 20468
rect 18844 20188 18900 20244
rect 18956 19964 19012 20020
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20748 23996 20804 24052
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 23212 28252 23268 28308
rect 22092 26962 22148 26964
rect 22092 26910 22094 26962
rect 22094 26910 22146 26962
rect 22146 26910 22148 26962
rect 22092 26908 22148 26910
rect 19964 23714 20020 23716
rect 19964 23662 19966 23714
rect 19966 23662 20018 23714
rect 20018 23662 20020 23714
rect 19964 23660 20020 23662
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19740 22258 19796 22260
rect 19740 22206 19742 22258
rect 19742 22206 19794 22258
rect 19794 22206 19796 22258
rect 19740 22204 19796 22206
rect 19964 22258 20020 22260
rect 19964 22206 19966 22258
rect 19966 22206 20018 22258
rect 20018 22206 20020 22258
rect 19964 22204 20020 22206
rect 19628 22092 19684 22148
rect 20188 22146 20244 22148
rect 20188 22094 20190 22146
rect 20190 22094 20242 22146
rect 20242 22094 20244 22146
rect 20188 22092 20244 22094
rect 19628 21868 19684 21924
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20412 22092 20468 22148
rect 20524 21756 20580 21812
rect 21532 23660 21588 23716
rect 21420 22988 21476 23044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 24556 28252 24612 28308
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 23212 26908 23268 26964
rect 22204 24892 22260 24948
rect 22428 26124 22484 26180
rect 25564 26402 25620 26404
rect 25564 26350 25566 26402
rect 25566 26350 25618 26402
rect 25618 26350 25620 26402
rect 25564 26348 25620 26350
rect 37884 26348 37940 26404
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 25788 24780 25844 24836
rect 22428 24668 22484 24724
rect 23772 24556 23828 24612
rect 22204 23884 22260 23940
rect 22092 23660 22148 23716
rect 21196 22146 21252 22148
rect 21196 22094 21198 22146
rect 21198 22094 21250 22146
rect 21250 22094 21252 22146
rect 21196 22092 21252 22094
rect 21532 21756 21588 21812
rect 19852 20690 19908 20692
rect 19852 20638 19854 20690
rect 19854 20638 19906 20690
rect 19906 20638 19908 20690
rect 19852 20636 19908 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20076 20188 20132 20244
rect 19740 20018 19796 20020
rect 19740 19966 19742 20018
rect 19742 19966 19794 20018
rect 19794 19966 19796 20018
rect 19740 19964 19796 19966
rect 19516 19852 19572 19908
rect 21532 20860 21588 20916
rect 21308 20802 21364 20804
rect 21308 20750 21310 20802
rect 21310 20750 21362 20802
rect 21362 20750 21364 20802
rect 21308 20748 21364 20750
rect 20188 20076 20244 20132
rect 20860 20130 20916 20132
rect 20860 20078 20862 20130
rect 20862 20078 20914 20130
rect 20914 20078 20916 20130
rect 20860 20076 20916 20078
rect 18956 18956 19012 19012
rect 19404 18844 19460 18900
rect 18956 18732 19012 18788
rect 18732 18620 18788 18676
rect 18508 18508 18564 18564
rect 19180 18674 19236 18676
rect 19180 18622 19182 18674
rect 19182 18622 19234 18674
rect 19234 18622 19236 18674
rect 19180 18620 19236 18622
rect 18396 18284 18452 18340
rect 18956 18284 19012 18340
rect 18844 18060 18900 18116
rect 17724 17388 17780 17444
rect 18956 17612 19012 17668
rect 18508 17052 18564 17108
rect 19068 17052 19124 17108
rect 19180 16940 19236 16996
rect 19964 19180 20020 19236
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19516 18508 19572 18564
rect 19628 18172 19684 18228
rect 19404 17666 19460 17668
rect 19404 17614 19406 17666
rect 19406 17614 19458 17666
rect 19458 17614 19460 17666
rect 19404 17612 19460 17614
rect 20076 18284 20132 18340
rect 20300 19292 20356 19348
rect 20412 19122 20468 19124
rect 20412 19070 20414 19122
rect 20414 19070 20466 19122
rect 20466 19070 20468 19122
rect 20412 19068 20468 19070
rect 20300 18956 20356 19012
rect 21196 19852 21252 19908
rect 20636 19292 20692 19348
rect 20748 18562 20804 18564
rect 20748 18510 20750 18562
rect 20750 18510 20802 18562
rect 20802 18510 20804 18562
rect 20748 18508 20804 18510
rect 21196 18508 21252 18564
rect 20636 18284 20692 18340
rect 20300 17890 20356 17892
rect 20300 17838 20302 17890
rect 20302 17838 20354 17890
rect 20354 17838 20356 17890
rect 20300 17836 20356 17838
rect 21420 18450 21476 18452
rect 21420 18398 21422 18450
rect 21422 18398 21474 18450
rect 21474 18398 21476 18450
rect 21420 18396 21476 18398
rect 21532 17836 21588 17892
rect 17724 15202 17780 15204
rect 17724 15150 17726 15202
rect 17726 15150 17778 15202
rect 17778 15150 17780 15202
rect 17724 15148 17780 15150
rect 15932 14530 15988 14532
rect 15932 14478 15934 14530
rect 15934 14478 15986 14530
rect 15986 14478 15988 14530
rect 15932 14476 15988 14478
rect 17388 14476 17444 14532
rect 18172 14252 18228 14308
rect 17388 13746 17444 13748
rect 17388 13694 17390 13746
rect 17390 13694 17442 13746
rect 17442 13694 17444 13746
rect 17388 13692 17444 13694
rect 18732 15372 18788 15428
rect 19180 15426 19236 15428
rect 19180 15374 19182 15426
rect 19182 15374 19234 15426
rect 19234 15374 19236 15426
rect 19180 15372 19236 15374
rect 19292 15202 19348 15204
rect 19292 15150 19294 15202
rect 19294 15150 19346 15202
rect 19346 15150 19348 15202
rect 19292 15148 19348 15150
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 21196 17052 21252 17108
rect 21532 17388 21588 17444
rect 21980 20300 22036 20356
rect 22764 23938 22820 23940
rect 22764 23886 22766 23938
rect 22766 23886 22818 23938
rect 22818 23886 22820 23938
rect 22764 23884 22820 23886
rect 23100 23826 23156 23828
rect 23100 23774 23102 23826
rect 23102 23774 23154 23826
rect 23154 23774 23156 23826
rect 23100 23772 23156 23774
rect 23996 23996 24052 24052
rect 24668 24722 24724 24724
rect 24668 24670 24670 24722
rect 24670 24670 24722 24722
rect 24722 24670 24724 24722
rect 24668 24668 24724 24670
rect 22316 23042 22372 23044
rect 22316 22990 22318 23042
rect 22318 22990 22370 23042
rect 22370 22990 22372 23042
rect 22316 22988 22372 22990
rect 22204 22204 22260 22260
rect 22540 22258 22596 22260
rect 22540 22206 22542 22258
rect 22542 22206 22594 22258
rect 22594 22206 22596 22258
rect 22540 22204 22596 22206
rect 23212 22092 23268 22148
rect 23884 22092 23940 22148
rect 24332 23884 24388 23940
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 25116 23938 25172 23940
rect 25116 23886 25118 23938
rect 25118 23886 25170 23938
rect 25170 23886 25172 23938
rect 25116 23884 25172 23886
rect 26572 25282 26628 25284
rect 26572 25230 26574 25282
rect 26574 25230 26626 25282
rect 26626 25230 26628 25282
rect 26572 25228 26628 25230
rect 39900 25564 39956 25620
rect 37660 25228 37716 25284
rect 40012 24892 40068 24948
rect 37660 24722 37716 24724
rect 37660 24670 37662 24722
rect 37662 24670 37714 24722
rect 37714 24670 37716 24722
rect 37660 24668 37716 24670
rect 26236 23884 26292 23940
rect 26348 24556 26404 24612
rect 25564 23772 25620 23828
rect 25340 23714 25396 23716
rect 25340 23662 25342 23714
rect 25342 23662 25394 23714
rect 25394 23662 25396 23714
rect 25340 23660 25396 23662
rect 24668 23548 24724 23604
rect 25228 23492 25284 23548
rect 22428 20524 22484 20580
rect 23100 20524 23156 20580
rect 22092 20076 22148 20132
rect 21980 18620 22036 18676
rect 21868 18562 21924 18564
rect 21868 18510 21870 18562
rect 21870 18510 21922 18562
rect 21922 18510 21924 18562
rect 21868 18508 21924 18510
rect 22428 18562 22484 18564
rect 22428 18510 22430 18562
rect 22430 18510 22482 18562
rect 22482 18510 22484 18562
rect 22428 18508 22484 18510
rect 21868 18226 21924 18228
rect 21868 18174 21870 18226
rect 21870 18174 21922 18226
rect 21922 18174 21924 18226
rect 21868 18172 21924 18174
rect 21756 17724 21812 17780
rect 21868 17836 21924 17892
rect 22540 18172 22596 18228
rect 24556 21420 24612 21476
rect 24220 21026 24276 21028
rect 24220 20974 24222 21026
rect 24222 20974 24274 21026
rect 24274 20974 24276 21026
rect 24220 20972 24276 20974
rect 24444 20914 24500 20916
rect 24444 20862 24446 20914
rect 24446 20862 24498 20914
rect 24498 20862 24500 20914
rect 24444 20860 24500 20862
rect 24668 20690 24724 20692
rect 24668 20638 24670 20690
rect 24670 20638 24722 20690
rect 24722 20638 24724 20690
rect 24668 20636 24724 20638
rect 24108 20524 24164 20580
rect 23996 20300 24052 20356
rect 28140 24610 28196 24612
rect 28140 24558 28142 24610
rect 28142 24558 28194 24610
rect 28194 24558 28196 24610
rect 28140 24556 28196 24558
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 40012 24220 40068 24276
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 26460 23826 26516 23828
rect 26460 23774 26462 23826
rect 26462 23774 26514 23826
rect 26514 23774 26516 23826
rect 26460 23772 26516 23774
rect 40012 23548 40068 23604
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 40012 22204 40068 22260
rect 37660 21756 37716 21812
rect 28812 21698 28868 21700
rect 28812 21646 28814 21698
rect 28814 21646 28866 21698
rect 28866 21646 28868 21698
rect 28812 21644 28868 21646
rect 28588 21586 28644 21588
rect 28588 21534 28590 21586
rect 28590 21534 28642 21586
rect 28642 21534 28644 21586
rect 28588 21532 28644 21534
rect 26012 21474 26068 21476
rect 26012 21422 26014 21474
rect 26014 21422 26066 21474
rect 26066 21422 26068 21474
rect 26012 21420 26068 21422
rect 27020 21420 27076 21476
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 40012 21532 40068 21588
rect 28140 21474 28196 21476
rect 28140 21422 28142 21474
rect 28142 21422 28194 21474
rect 28194 21422 28196 21474
rect 28140 21420 28196 21422
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 26908 20690 26964 20692
rect 26908 20638 26910 20690
rect 26910 20638 26962 20690
rect 26962 20638 26964 20690
rect 26908 20636 26964 20638
rect 25452 20188 25508 20244
rect 25900 20300 25956 20356
rect 23772 19628 23828 19684
rect 23436 18396 23492 18452
rect 23772 19068 23828 19124
rect 24220 19068 24276 19124
rect 21756 16828 21812 16884
rect 23212 16098 23268 16100
rect 23212 16046 23214 16098
rect 23214 16046 23266 16098
rect 23266 16046 23268 16098
rect 23212 16044 23268 16046
rect 25228 19628 25284 19684
rect 25116 19234 25172 19236
rect 25116 19182 25118 19234
rect 25118 19182 25170 19234
rect 25170 19182 25172 19234
rect 25116 19180 25172 19182
rect 25788 19852 25844 19908
rect 25564 19122 25620 19124
rect 25564 19070 25566 19122
rect 25566 19070 25618 19122
rect 25618 19070 25620 19122
rect 25564 19068 25620 19070
rect 28364 19906 28420 19908
rect 28364 19854 28366 19906
rect 28366 19854 28418 19906
rect 28418 19854 28420 19906
rect 28364 19852 28420 19854
rect 40012 20188 40068 20244
rect 37660 19852 37716 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 26348 19068 26404 19124
rect 25340 18396 25396 18452
rect 25676 18450 25732 18452
rect 25676 18398 25678 18450
rect 25678 18398 25730 18450
rect 25730 18398 25732 18450
rect 25676 18396 25732 18398
rect 26124 18450 26180 18452
rect 26124 18398 26126 18450
rect 26126 18398 26178 18450
rect 26178 18398 26180 18450
rect 26124 18396 26180 18398
rect 25452 18338 25508 18340
rect 25452 18286 25454 18338
rect 25454 18286 25506 18338
rect 25506 18286 25508 18338
rect 25452 18284 25508 18286
rect 24332 16828 24388 16884
rect 25228 17106 25284 17108
rect 25228 17054 25230 17106
rect 25230 17054 25282 17106
rect 25282 17054 25284 17106
rect 25228 17052 25284 17054
rect 26236 16994 26292 16996
rect 26236 16942 26238 16994
rect 26238 16942 26290 16994
rect 26290 16942 26292 16994
rect 26236 16940 26292 16942
rect 27020 18396 27076 18452
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 27132 17052 27188 17108
rect 21532 15372 21588 15428
rect 21196 15314 21252 15316
rect 21196 15262 21198 15314
rect 21198 15262 21250 15314
rect 21250 15262 21252 15314
rect 21196 15260 21252 15262
rect 19964 15148 20020 15204
rect 18732 14588 18788 14644
rect 19516 14642 19572 14644
rect 19516 14590 19518 14642
rect 19518 14590 19570 14642
rect 19570 14590 19572 14642
rect 19516 14588 19572 14590
rect 18620 13692 18676 13748
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 21644 15148 21700 15204
rect 20748 14588 20804 14644
rect 19852 14306 19908 14308
rect 19852 14254 19854 14306
rect 19854 14254 19906 14306
rect 19906 14254 19908 14306
rect 19852 14252 19908 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 23884 16098 23940 16100
rect 23884 16046 23886 16098
rect 23886 16046 23938 16098
rect 23938 16046 23940 16098
rect 23884 16044 23940 16046
rect 28028 17052 28084 17108
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37660 17052 37716 17108
rect 27580 16828 27636 16884
rect 37660 16882 37716 16884
rect 37660 16830 37662 16882
rect 37662 16830 37714 16882
rect 37714 16830 37716 16882
rect 37660 16828 37716 16830
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 40012 16156 40068 16212
rect 26348 16044 26404 16100
rect 23660 15874 23716 15876
rect 23660 15822 23662 15874
rect 23662 15822 23714 15874
rect 23714 15822 23716 15874
rect 23660 15820 23716 15822
rect 25788 15820 25844 15876
rect 23436 15260 23492 15316
rect 22092 14642 22148 14644
rect 22092 14590 22094 14642
rect 22094 14590 22146 14642
rect 22146 14590 22148 14642
rect 22092 14588 22148 14590
rect 22876 14588 22932 14644
rect 23996 14588 24052 14644
rect 20748 13746 20804 13748
rect 20748 13694 20750 13746
rect 20750 13694 20802 13746
rect 20802 13694 20804 13746
rect 20748 13692 20804 13694
rect 19628 13132 19684 13188
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 22540 13468 22596 13524
rect 23548 13468 23604 13524
rect 24556 13468 24612 13524
rect 20636 13186 20692 13188
rect 20636 13134 20638 13186
rect 20638 13134 20690 13186
rect 20690 13134 20692 13186
rect 20636 13132 20692 13134
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18844 4060 18900 4116
rect 20076 4114 20132 4116
rect 20076 4062 20078 4114
rect 20078 4062 20130 4114
rect 20130 4062 20132 4114
rect 20076 4060 20132 4062
rect 20860 3612 20916 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 24220 4060 24276 4116
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 22876 3612 22932 3668
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 14914 37996 14924 38052
rect 14980 37996 15932 38052
rect 15988 37996 15998 38052
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16146 37436 16156 37492
rect 16212 37436 18396 37492
rect 18452 37436 18462 37492
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 0 37044 800 37072
rect 0 36988 1708 37044
rect 1764 36988 1774 37044
rect 0 36960 800 36988
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 15474 36652 15484 36708
rect 15540 36652 16716 36708
rect 16772 36652 16782 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 14578 28588 14588 28644
rect 14644 28588 16268 28644
rect 16324 28588 16828 28644
rect 16884 28588 16894 28644
rect 13458 28476 13468 28532
rect 13524 28476 14924 28532
rect 14980 28476 14990 28532
rect 17378 28476 17388 28532
rect 17444 28476 18620 28532
rect 18676 28476 18686 28532
rect 0 28308 800 28336
rect 0 28252 4172 28308
rect 4228 28252 4238 28308
rect 23202 28252 23212 28308
rect 23268 28252 24556 28308
rect 24612 28252 24622 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 14354 27468 14364 27524
rect 14420 27468 15708 27524
rect 15764 27468 15774 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 1922 27132 1932 27188
rect 1988 27132 1998 27188
rect 13906 27132 13916 27188
rect 13972 27132 15148 27188
rect 15204 27132 15876 27188
rect 0 26964 800 26992
rect 1932 26964 1988 27132
rect 15820 27076 15876 27132
rect 4274 27020 4284 27076
rect 4340 27020 11228 27076
rect 11284 27020 13804 27076
rect 13860 27020 13870 27076
rect 14914 27020 14924 27076
rect 14980 27020 15596 27076
rect 15652 27020 15662 27076
rect 15810 27020 15820 27076
rect 15876 27020 17948 27076
rect 18004 27020 18014 27076
rect 0 26908 1988 26964
rect 13122 26908 13132 26964
rect 13188 26908 14252 26964
rect 14308 26908 14318 26964
rect 15026 26908 15036 26964
rect 15092 26908 17276 26964
rect 17332 26908 17342 26964
rect 22082 26908 22092 26964
rect 22148 26908 23212 26964
rect 23268 26908 23278 26964
rect 0 26880 800 26908
rect 14466 26796 14476 26852
rect 14532 26796 15372 26852
rect 15428 26796 15438 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 25554 26348 25564 26404
rect 25620 26348 37884 26404
rect 37940 26348 37950 26404
rect 14130 26124 14140 26180
rect 14196 26124 15708 26180
rect 15764 26124 17724 26180
rect 17780 26124 19516 26180
rect 19572 26124 19964 26180
rect 20020 26124 20412 26180
rect 20468 26124 22428 26180
rect 22484 26124 22494 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 13346 25676 13356 25732
rect 13412 25676 13916 25732
rect 13972 25676 13982 25732
rect 41200 25620 42000 25648
rect 39890 25564 39900 25620
rect 39956 25564 42000 25620
rect 41200 25536 42000 25564
rect 12450 25228 12460 25284
rect 12516 25228 14084 25284
rect 26562 25228 26572 25284
rect 26628 25228 37660 25284
rect 37716 25228 37726 25284
rect 14028 25060 14084 25228
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 14018 25004 14028 25060
rect 14084 25004 14094 25060
rect 41200 24948 42000 24976
rect 13458 24892 13468 24948
rect 13524 24892 15148 24948
rect 15204 24892 15214 24948
rect 18162 24892 18172 24948
rect 18228 24892 22204 24948
rect 22260 24892 22270 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 41200 24864 42000 24892
rect 17490 24780 17500 24836
rect 17556 24780 18284 24836
rect 18340 24780 19292 24836
rect 19348 24780 19358 24836
rect 25778 24780 25788 24836
rect 25844 24780 25854 24836
rect 22418 24668 22428 24724
rect 22484 24668 24668 24724
rect 24724 24668 25228 24724
rect 25284 24668 25294 24724
rect 25788 24612 25844 24780
rect 31892 24668 37660 24724
rect 37716 24668 37726 24724
rect 31892 24612 31948 24668
rect 23762 24556 23772 24612
rect 23828 24556 25844 24612
rect 26338 24556 26348 24612
rect 26404 24556 28140 24612
rect 28196 24556 31948 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 20524 23996 20748 24052
rect 20804 23996 23996 24052
rect 24052 23996 24062 24052
rect 13794 23884 13804 23940
rect 13860 23884 14588 23940
rect 14644 23884 14654 23940
rect 20524 23828 20580 23996
rect 22194 23884 22204 23940
rect 22260 23884 22764 23940
rect 22820 23884 22830 23940
rect 24322 23884 24332 23940
rect 24388 23884 25116 23940
rect 25172 23884 25182 23940
rect 26226 23884 26236 23940
rect 26292 23884 37660 23940
rect 37716 23884 37726 23940
rect 14354 23772 14364 23828
rect 14420 23772 15036 23828
rect 15092 23772 17836 23828
rect 17892 23772 17902 23828
rect 19394 23772 19404 23828
rect 19460 23772 20580 23828
rect 23090 23772 23100 23828
rect 23156 23772 25564 23828
rect 25620 23772 26460 23828
rect 26516 23772 26526 23828
rect 13682 23660 13692 23716
rect 13748 23660 14140 23716
rect 14196 23660 14206 23716
rect 15138 23660 15148 23716
rect 15204 23660 17500 23716
rect 17556 23660 19964 23716
rect 20020 23660 21532 23716
rect 21588 23660 21598 23716
rect 22082 23660 22092 23716
rect 22148 23660 25340 23716
rect 25396 23660 25406 23716
rect 41200 23604 42000 23632
rect 24658 23548 24668 23604
rect 24724 23548 25284 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 25218 23492 25228 23548
rect 25284 23492 25294 23548
rect 41200 23520 42000 23548
rect 15138 23212 15148 23268
rect 15204 23212 15820 23268
rect 15876 23212 15886 23268
rect 11666 22988 11676 23044
rect 11732 22988 14252 23044
rect 14308 22988 14318 23044
rect 17490 22988 17500 23044
rect 17556 22988 18172 23044
rect 18228 22988 18238 23044
rect 21410 22988 21420 23044
rect 21476 22988 22316 23044
rect 22372 22988 22382 23044
rect 13906 22876 13916 22932
rect 13972 22876 14924 22932
rect 14980 22876 14990 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 16146 22316 16156 22372
rect 16212 22316 17612 22372
rect 17668 22316 17678 22372
rect 41200 22260 42000 22288
rect 14578 22204 14588 22260
rect 14644 22204 15932 22260
rect 15988 22204 15998 22260
rect 17154 22204 17164 22260
rect 17220 22204 17388 22260
rect 17444 22204 17454 22260
rect 18498 22204 18508 22260
rect 18564 22204 19740 22260
rect 19796 22204 19806 22260
rect 19954 22204 19964 22260
rect 20020 22204 22204 22260
rect 22260 22204 22540 22260
rect 22596 22204 22606 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 4162 22092 4172 22148
rect 4228 22092 18620 22148
rect 18676 22092 18686 22148
rect 19618 22092 19628 22148
rect 19684 22092 20188 22148
rect 20244 22092 20254 22148
rect 20402 22092 20412 22148
rect 20468 22092 21196 22148
rect 21252 22092 21262 22148
rect 23202 22092 23212 22148
rect 23268 22092 23884 22148
rect 23940 22092 23950 22148
rect 10994 21980 11004 22036
rect 11060 21980 13132 22036
rect 13188 21980 14028 22036
rect 14084 21980 14094 22036
rect 14466 21980 14476 22036
rect 14532 21980 17164 22036
rect 17220 21980 17230 22036
rect 17490 21980 17500 22036
rect 17556 21980 19292 22036
rect 19348 21980 19358 22036
rect 14476 21924 14532 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 13906 21868 13916 21924
rect 13972 21868 14532 21924
rect 15810 21868 15820 21924
rect 15876 21868 19628 21924
rect 19684 21868 19694 21924
rect 14018 21644 14028 21700
rect 14084 21644 14476 21700
rect 14532 21644 14924 21700
rect 14980 21644 14990 21700
rect 4274 21532 4284 21588
rect 4340 21532 9996 21588
rect 10052 21532 10062 21588
rect 17724 21476 17780 21868
rect 20514 21756 20524 21812
rect 20580 21756 21532 21812
rect 21588 21756 21598 21812
rect 31892 21756 37660 21812
rect 37716 21756 37726 21812
rect 31892 21700 31948 21756
rect 28802 21644 28812 21700
rect 28868 21644 31948 21700
rect 41200 21588 42000 21616
rect 28578 21532 28588 21588
rect 28644 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 17714 21420 17724 21476
rect 17780 21420 17790 21476
rect 24546 21420 24556 21476
rect 24612 21420 26012 21476
rect 26068 21420 26078 21476
rect 27010 21420 27020 21476
rect 27076 21420 28140 21476
rect 28196 21420 28206 21476
rect 17490 21308 17500 21364
rect 17556 21308 18172 21364
rect 18228 21308 18620 21364
rect 18676 21308 18686 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 17938 20972 17948 21028
rect 18004 20972 24220 21028
rect 24276 20972 24286 21028
rect 0 20916 800 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 9986 20860 9996 20916
rect 10052 20860 14700 20916
rect 14756 20860 14766 20916
rect 16370 20860 16380 20916
rect 16436 20860 17164 20916
rect 17220 20860 17230 20916
rect 21522 20860 21532 20916
rect 21588 20860 24444 20916
rect 24500 20860 24510 20916
rect 0 20832 800 20860
rect 13570 20748 13580 20804
rect 13636 20748 15708 20804
rect 15764 20748 15774 20804
rect 16146 20748 16156 20804
rect 16212 20748 17388 20804
rect 17444 20748 17454 20804
rect 18498 20748 18508 20804
rect 18564 20748 21308 20804
rect 21364 20748 21374 20804
rect 12114 20636 12124 20692
rect 12180 20636 15372 20692
rect 15428 20636 15438 20692
rect 18722 20636 18732 20692
rect 18788 20636 19852 20692
rect 19908 20636 19918 20692
rect 24658 20636 24668 20692
rect 24724 20636 26908 20692
rect 26964 20636 26974 20692
rect 12226 20524 12236 20580
rect 12292 20524 13804 20580
rect 13860 20524 13870 20580
rect 19180 20524 22428 20580
rect 22484 20524 23100 20580
rect 23156 20524 24108 20580
rect 24164 20524 24174 20580
rect 19180 20468 19236 20524
rect 14802 20412 14812 20468
rect 14868 20412 19180 20468
rect 19236 20412 19246 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 21970 20300 21980 20356
rect 22036 20300 23996 20356
rect 24052 20300 25900 20356
rect 25956 20300 25966 20356
rect 41200 20244 42000 20272
rect 17714 20188 17724 20244
rect 17780 20188 18844 20244
rect 18900 20188 20076 20244
rect 20132 20188 20142 20244
rect 25442 20188 25452 20244
rect 25508 20188 25564 20244
rect 25620 20188 25630 20244
rect 40002 20188 40012 20244
rect 40068 20188 42000 20244
rect 41200 20160 42000 20188
rect 15250 20076 15260 20132
rect 15316 20076 18060 20132
rect 18116 20076 18126 20132
rect 18834 20076 18844 20132
rect 18900 20076 20188 20132
rect 20244 20076 20254 20132
rect 20850 20076 20860 20132
rect 20916 20076 22092 20132
rect 22148 20076 22158 20132
rect 18946 19964 18956 20020
rect 19012 19964 19740 20020
rect 19796 19964 19806 20020
rect 19506 19852 19516 19908
rect 19572 19852 21196 19908
rect 21252 19852 21262 19908
rect 25778 19852 25788 19908
rect 25844 19852 28364 19908
rect 28420 19852 37660 19908
rect 37716 19852 37726 19908
rect 23762 19628 23772 19684
rect 23828 19628 25228 19684
rect 25284 19628 25294 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 14354 19404 14364 19460
rect 14420 19404 14924 19460
rect 14980 19404 15148 19460
rect 15474 19404 15484 19460
rect 15540 19404 20356 19460
rect 15092 19348 15148 19404
rect 20300 19348 20356 19404
rect 15092 19292 17836 19348
rect 17892 19292 17902 19348
rect 20290 19292 20300 19348
rect 20356 19292 20636 19348
rect 20692 19292 20702 19348
rect 14242 19180 14252 19236
rect 14308 19180 14924 19236
rect 14980 19180 16156 19236
rect 16212 19180 17052 19236
rect 17108 19180 17118 19236
rect 18050 19180 18060 19236
rect 18116 19180 19964 19236
rect 20020 19180 25116 19236
rect 25172 19180 25182 19236
rect 16370 19068 16380 19124
rect 16436 19068 20412 19124
rect 20468 19068 23772 19124
rect 23828 19068 24220 19124
rect 24276 19068 24286 19124
rect 25526 19068 25564 19124
rect 25620 19068 26348 19124
rect 26404 19068 26414 19124
rect 18050 18956 18060 19012
rect 18116 18956 18956 19012
rect 19012 18956 19022 19012
rect 19404 18956 20300 19012
rect 20356 18956 20366 19012
rect 19404 18900 19460 18956
rect 17378 18844 17388 18900
rect 17444 18844 19404 18900
rect 19460 18844 19470 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 16818 18732 16828 18788
rect 16884 18732 18284 18788
rect 18340 18732 18956 18788
rect 19012 18732 19022 18788
rect 18722 18620 18732 18676
rect 18788 18620 19180 18676
rect 19236 18620 19246 18676
rect 21634 18620 21644 18676
rect 21700 18620 21980 18676
rect 22036 18620 22046 18676
rect 18498 18508 18508 18564
rect 18564 18508 19516 18564
rect 19572 18508 19582 18564
rect 20738 18508 20748 18564
rect 20804 18508 21196 18564
rect 21252 18508 21868 18564
rect 21924 18508 22428 18564
rect 22484 18508 22494 18564
rect 11442 18396 11452 18452
rect 11508 18396 15036 18452
rect 15092 18396 15102 18452
rect 17938 18396 17948 18452
rect 18004 18396 21420 18452
rect 21476 18396 21486 18452
rect 23426 18396 23436 18452
rect 23492 18396 25340 18452
rect 25396 18396 25676 18452
rect 25732 18396 25742 18452
rect 26114 18396 26124 18452
rect 26180 18396 27020 18452
rect 27076 18396 27086 18452
rect 14914 18284 14924 18340
rect 14980 18284 16492 18340
rect 16548 18284 17052 18340
rect 17108 18284 17118 18340
rect 17714 18284 17724 18340
rect 17780 18284 18396 18340
rect 18452 18284 18956 18340
rect 19012 18284 19022 18340
rect 20066 18284 20076 18340
rect 20132 18284 20636 18340
rect 20692 18284 25452 18340
rect 25508 18284 25518 18340
rect 41200 18228 42000 18256
rect 19618 18172 19628 18228
rect 19684 18172 21868 18228
rect 21924 18172 22540 18228
rect 22596 18172 22606 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 18806 18060 18844 18116
rect 18900 18060 18910 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 15474 17836 15484 17892
rect 15540 17836 17948 17892
rect 18004 17836 18014 17892
rect 20290 17836 20300 17892
rect 20356 17836 21532 17892
rect 21588 17836 21868 17892
rect 21924 17836 21934 17892
rect 21532 17724 21756 17780
rect 21812 17724 21822 17780
rect 4274 17612 4284 17668
rect 4340 17612 12012 17668
rect 12068 17612 15260 17668
rect 15316 17612 15326 17668
rect 17378 17612 17388 17668
rect 17444 17612 18956 17668
rect 19012 17612 19404 17668
rect 19460 17612 19470 17668
rect 21532 17444 21588 17724
rect 14914 17388 14924 17444
rect 14980 17388 15484 17444
rect 15540 17388 17724 17444
rect 17780 17388 17790 17444
rect 21522 17388 21532 17444
rect 21588 17388 21598 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 11788 17052 15372 17108
rect 15428 17052 15438 17108
rect 18498 17052 18508 17108
rect 18564 17052 19068 17108
rect 19124 17052 21196 17108
rect 21252 17052 25228 17108
rect 25284 17052 25294 17108
rect 27122 17052 27132 17108
rect 27188 17052 28028 17108
rect 28084 17052 37660 17108
rect 37716 17052 37726 17108
rect 11788 16996 11844 17052
rect 4274 16940 4284 16996
rect 4340 16940 11788 16996
rect 11844 16940 11854 16996
rect 14802 16940 14812 16996
rect 14868 16940 19180 16996
rect 19236 16940 19246 16996
rect 26226 16940 26236 16996
rect 26292 16940 26908 16996
rect 0 16884 800 16912
rect 26852 16884 26908 16940
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 14466 16828 14476 16884
rect 14532 16828 15372 16884
rect 15428 16828 15438 16884
rect 21746 16828 21756 16884
rect 21812 16828 24332 16884
rect 24388 16828 24398 16884
rect 26852 16828 27580 16884
rect 27636 16828 37660 16884
rect 37716 16828 37726 16884
rect 0 16800 800 16828
rect 15138 16716 15148 16772
rect 15204 16716 15932 16772
rect 15988 16716 15998 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16212 800 16240
rect 41200 16212 42000 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 40002 16156 40012 16212
rect 40068 16156 42000 16212
rect 0 16128 800 16156
rect 41200 16128 42000 16156
rect 14242 16044 14252 16100
rect 14308 16044 23212 16100
rect 23268 16044 23278 16100
rect 23874 16044 23884 16100
rect 23940 16044 26348 16100
rect 26404 16044 26414 16100
rect 23650 15820 23660 15876
rect 23716 15820 25788 15876
rect 25844 15820 25854 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 18722 15372 18732 15428
rect 18788 15372 19180 15428
rect 19236 15372 21532 15428
rect 21588 15372 21598 15428
rect 21186 15260 21196 15316
rect 21252 15260 23436 15316
rect 23492 15260 23502 15316
rect 17714 15148 17724 15204
rect 17780 15148 19292 15204
rect 19348 15148 19358 15204
rect 19954 15148 19964 15204
rect 20020 15148 21644 15204
rect 21700 15148 21710 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 18722 14588 18732 14644
rect 18788 14588 19516 14644
rect 19572 14588 19582 14644
rect 20738 14588 20748 14644
rect 20804 14588 22092 14644
rect 22148 14588 22876 14644
rect 22932 14588 23996 14644
rect 24052 14588 24062 14644
rect 15922 14476 15932 14532
rect 15988 14476 17388 14532
rect 17444 14476 17454 14532
rect 18162 14252 18172 14308
rect 18228 14252 19852 14308
rect 19908 14252 19918 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 17378 13692 17388 13748
rect 17444 13692 18620 13748
rect 18676 13692 20748 13748
rect 20804 13692 20814 13748
rect 22530 13468 22540 13524
rect 22596 13468 23548 13524
rect 23604 13468 24556 13524
rect 24612 13468 24622 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19618 13132 19628 13188
rect 19684 13132 20636 13188
rect 20692 13132 20702 13188
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 18834 4060 18844 4116
rect 18900 4060 20076 4116
rect 20132 4060 20142 4116
rect 24210 4060 24220 4116
rect 24276 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 22866 3612 22876 3668
rect 22932 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 25564 20188 25620 20244
rect 18844 20076 18900 20132
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 25564 19068 25620 19124
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 21644 18620 21700 18676
rect 18844 18060 18900 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 21644 15148 21700 15204
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 18844 20132 18900 20142
rect 18844 18116 18900 20076
rect 18844 18050 18900 18060
rect 19808 18844 20128 20356
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 25564 20244 25620 20254
rect 25564 19124 25620 20188
rect 25564 19058 25620 19068
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 21644 18676 21700 18686
rect 21644 15204 21700 18620
rect 21644 15138 21700 15148
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24080 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform 1 0 18480 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14784 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18592 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform 1 0 22624 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 25984 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _107_
timestamp 1698175906
transform 1 0 25872 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform 1 0 20272 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _109_
timestamp 1698175906
transform -1 0 22624 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14784 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19600 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform 1 0 17024 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14672 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 20048 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _116_
timestamp 1698175906
transform -1 0 19824 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform 1 0 18032 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _122_
timestamp 1698175906
transform -1 0 17920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform 1 0 18704 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 23856 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21728 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform -1 0 26544 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _128_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16576 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform -1 0 16352 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16688 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _132_
timestamp 1698175906
transform -1 0 14112 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _133_
timestamp 1698175906
transform 1 0 15680 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 14448 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14896 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform 1 0 14000 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _137_
timestamp 1698175906
transform 1 0 17808 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 15904 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _139_
timestamp 1698175906
transform 1 0 14784 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_
timestamp 1698175906
transform 1 0 19488 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform 1 0 22288 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _142_
timestamp 1698175906
transform 1 0 22960 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _143_
timestamp 1698175906
transform 1 0 23296 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform 1 0 23520 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform -1 0 18480 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 15344 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _147_
timestamp 1698175906
transform -1 0 14784 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _148_
timestamp 1698175906
transform 1 0 21728 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _149_
timestamp 1698175906
transform -1 0 22176 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform -1 0 26656 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _151_
timestamp 1698175906
transform 1 0 24976 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _152_
timestamp 1698175906
transform -1 0 22512 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _153_
timestamp 1698175906
transform -1 0 27328 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18704 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _156_
timestamp 1698175906
transform 1 0 19936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform 1 0 20944 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform 1 0 18368 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 18928 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform -1 0 18256 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _161_
timestamp 1698175906
transform -1 0 18928 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 21728 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _163_
timestamp 1698175906
transform -1 0 20496 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _164_
timestamp 1698175906
transform -1 0 18480 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1698175906
transform 1 0 17584 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _166_
timestamp 1698175906
transform 1 0 14784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform -1 0 14784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform 1 0 22512 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698175906
transform -1 0 22736 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _170_
timestamp 1698175906
transform 1 0 20832 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform -1 0 15680 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform -1 0 14896 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform -1 0 15008 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14448 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _176_
timestamp 1698175906
transform -1 0 27216 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _177_
timestamp 1698175906
transform 1 0 23632 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _178_
timestamp 1698175906
transform 1 0 23072 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _179_
timestamp 1698175906
transform -1 0 24080 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform -1 0 19264 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _182_
timestamp 1698175906
transform -1 0 17024 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform -1 0 14784 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform -1 0 15904 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform -1 0 16016 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform 1 0 13216 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform -1 0 14112 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _188_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13664 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _189_
timestamp 1698175906
transform -1 0 20944 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698175906
transform 1 0 17248 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 22400 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _193_
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 17584 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 15792 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform 1 0 24528 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 10752 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 13776 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22624 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 12208 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 24976 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform -1 0 20496 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 19264 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform -1 0 15120 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 20496 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform -1 0 14896 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform -1 0 13104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 22736 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 15008 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform -1 0 16576 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform -1 0 14336 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 20160 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _220_
timestamp 1698175906
transform 1 0 28336 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _221_
timestamp 1698175906
transform 1 0 26096 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _222_
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _223_
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 19936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform -1 0 19264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 24304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform -1 0 21504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform -1 0 15456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 14000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 22400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 15680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 24752 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 20720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 22736 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 15904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 23968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform -1 0 18704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 16800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 19488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18256 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 24528 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform -1 0 23520 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 23632 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_115
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_119
timestamp 1698175906
transform 1 0 14672 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_121
timestamp 1698175906
transform 1 0 14896 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_151
timestamp 1698175906
transform 1 0 18256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_155
timestamp 1698175906
transform 1 0 18704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_157
timestamp 1698175906
transform 1 0 18928 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_160
timestamp 1698175906
transform 1 0 19264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_168
timestamp 1698175906
transform 1 0 20160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_170
timestamp 1698175906
transform 1 0 20384 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_200
timestamp 1698175906
transform 1 0 23744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_204
timestamp 1698175906
transform 1 0 24192 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_127
timestamp 1698175906
transform 1 0 15568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_158
timestamp 1698175906
transform 1 0 19040 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_169
timestamp 1698175906
transform 1 0 20272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_220
timestamp 1698175906
transform 1 0 25984 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_236
timestamp 1698175906
transform 1 0 27776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_121
timestamp 1698175906
transform 1 0 14896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_125
timestamp 1698175906
transform 1 0 15344 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698175906
transform 1 0 16240 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698175906
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_166
timestamp 1698175906
transform 1 0 19936 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_186
timestamp 1698175906
transform 1 0 22176 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_194
timestamp 1698175906
transform 1 0 23072 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_198
timestamp 1698175906
transform 1 0 23520 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698175906
transform 1 0 24080 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698175906
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_121
timestamp 1698175906
transform 1 0 14896 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_153
timestamp 1698175906
transform 1 0 18480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_160
timestamp 1698175906
transform 1 0 19264 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1698175906
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_193
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_203
timestamp 1698175906
transform 1 0 24080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_236
timestamp 1698175906
transform 1 0 27776 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_92
timestamp 1698175906
transform 1 0 11648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_128
timestamp 1698175906
transform 1 0 15680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_132
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698175906
transform 1 0 18144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_154
timestamp 1698175906
transform 1 0 18592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_156
timestamp 1698175906
transform 1 0 18816 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_225
timestamp 1698175906
transform 1 0 26544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_227
timestamp 1698175906
transform 1 0 26768 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_232
timestamp 1698175906
transform 1 0 27328 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_264
timestamp 1698175906
transform 1 0 30912 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_128
timestamp 1698175906
transform 1 0 15680 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_136
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_138
timestamp 1698175906
transform 1 0 16800 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_145
timestamp 1698175906
transform 1 0 17584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_186
timestamp 1698175906
transform 1 0 22176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_188
timestamp 1698175906
transform 1 0 22400 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_195
timestamp 1698175906
transform 1 0 23184 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_203
timestamp 1698175906
transform 1 0 24080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_207
timestamp 1698175906
transform 1 0 24528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 28224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_120
timestamp 1698175906
transform 1 0 14784 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_128
timestamp 1698175906
transform 1 0 15680 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_132
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_190
timestamp 1698175906
transform 1 0 22624 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_194
timestamp 1698175906
transform 1 0 23072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_196
timestamp 1698175906
transform 1 0 23296 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_224
timestamp 1698175906
transform 1 0 26432 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_256
timestamp 1698175906
transform 1 0 30016 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_272
timestamp 1698175906
transform 1 0 31808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_136
timestamp 1698175906
transform 1 0 16576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_138
timestamp 1698175906
transform 1 0 16800 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_151
timestamp 1698175906
transform 1 0 18256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_153
timestamp 1698175906
transform 1 0 18480 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_168
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_206
timestamp 1698175906
transform 1 0 24416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_210
timestamp 1698175906
transform 1 0 24864 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_220
timestamp 1698175906
transform 1 0 25984 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_236
timestamp 1698175906
transform 1 0 27776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_122
timestamp 1698175906
transform 1 0 15008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_126
timestamp 1698175906
transform 1 0 15456 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_146
timestamp 1698175906
transform 1 0 17696 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_159
timestamp 1698175906
transform 1 0 19152 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_176
timestamp 1698175906
transform 1 0 21056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_180
timestamp 1698175906
transform 1 0 21504 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_196
timestamp 1698175906
transform 1 0 23296 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_204
timestamp 1698175906
transform 1 0 24192 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_243
timestamp 1698175906
transform 1 0 28560 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698175906
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 9744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_114
timestamp 1698175906
transform 1 0 14112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_116
timestamp 1698175906
transform 1 0 14336 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_134
timestamp 1698175906
transform 1 0 16352 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_138
timestamp 1698175906
transform 1 0 16800 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_153
timestamp 1698175906
transform 1 0 18480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_161
timestamp 1698175906
transform 1 0 19376 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_189
timestamp 1698175906
transform 1 0 22512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_210
timestamp 1698175906
transform 1 0 24864 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_218
timestamp 1698175906
transform 1 0 25760 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_223
timestamp 1698175906
transform 1 0 26320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_231
timestamp 1698175906
transform 1 0 27216 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_239
timestamp 1698175906
transform 1 0 28112 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698175906
transform 1 0 12992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_107
timestamp 1698175906
transform 1 0 13328 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_115
timestamp 1698175906
transform 1 0 14224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_123
timestamp 1698175906
transform 1 0 15120 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_247
timestamp 1698175906
transform 1 0 29008 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_124
timestamp 1698175906
transform 1 0 15232 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_134
timestamp 1698175906
transform 1 0 16352 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_148
timestamp 1698175906
transform 1 0 17920 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_155
timestamp 1698175906
transform 1 0 18704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_159
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_161
timestamp 1698175906
transform 1 0 19376 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698175906
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_182
timestamp 1698175906
transform 1 0 21728 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_186
timestamp 1698175906
transform 1 0 22176 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_192
timestamp 1698175906
transform 1 0 22848 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_208
timestamp 1698175906
transform 1 0 24640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_212
timestamp 1698175906
transform 1 0 25088 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_130
timestamp 1698175906
transform 1 0 15904 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_147
timestamp 1698175906
transform 1 0 17808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_155
timestamp 1698175906
transform 1 0 18704 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_159
timestamp 1698175906
transform 1 0 19152 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_189
timestamp 1698175906
transform 1 0 22512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_193
timestamp 1698175906
transform 1 0 22960 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_121
timestamp 1698175906
transform 1 0 14896 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_137
timestamp 1698175906
transform 1 0 16688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_139
timestamp 1698175906
transform 1 0 16912 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_152
timestamp 1698175906
transform 1 0 18368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_156
timestamp 1698175906
transform 1 0 18816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_158
timestamp 1698175906
transform 1 0 19040 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_173
timestamp 1698175906
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698175906
transform 1 0 22288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_204
timestamp 1698175906
transform 1 0 24192 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_208
timestamp 1698175906
transform 1 0 24640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_210
timestamp 1698175906
transform 1 0 24864 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_219
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_226
timestamp 1698175906
transform 1 0 26656 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_104
timestamp 1698175906
transform 1 0 12992 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_146
timestamp 1698175906
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698175906
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_241
timestamp 1698175906
transform 1 0 28336 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 31920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698175906
transform 1 0 13552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_117
timestamp 1698175906
transform 1 0 14448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_119
timestamp 1698175906
transform 1 0 14672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_128
timestamp 1698175906
transform 1 0 15680 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_144
timestamp 1698175906
transform 1 0 17472 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_188
timestamp 1698175906
transform 1 0 22400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_227
timestamp 1698175906
transform 1 0 26768 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_96
timestamp 1698175906
transform 1 0 12096 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_126
timestamp 1698175906
transform 1 0 15456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_130
timestamp 1698175906
transform 1 0 15904 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_153
timestamp 1698175906
transform 1 0 18480 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_161
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_164
timestamp 1698175906
transform 1 0 19712 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_197
timestamp 1698175906
transform 1 0 23408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698175906
transform 1 0 24304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_218
timestamp 1698175906
transform 1 0 25760 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_250
timestamp 1698175906
transform 1 0 29344 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_266
timestamp 1698175906
transform 1 0 31136 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698175906
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_114
timestamp 1698175906
transform 1 0 14112 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_130
timestamp 1698175906
transform 1 0 15904 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_146
timestamp 1698175906
transform 1 0 17696 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_154
timestamp 1698175906
transform 1 0 18592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_156
timestamp 1698175906
transform 1 0 18816 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_162
timestamp 1698175906
transform 1 0 19488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_170
timestamp 1698175906
transform 1 0 20384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698175906
transform 1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_188
timestamp 1698175906
transform 1 0 22400 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_220
timestamp 1698175906
transform 1 0 25984 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_236
timestamp 1698175906
transform 1 0 27776 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_80
timestamp 1698175906
transform 1 0 10304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_84
timestamp 1698175906
transform 1 0 10752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_86
timestamp 1698175906
transform 1 0 10976 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_116
timestamp 1698175906
transform 1 0 14336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_131
timestamp 1698175906
transform 1 0 16016 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_171
timestamp 1698175906
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_175
timestamp 1698175906
transform 1 0 20944 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_136
timestamp 1698175906
transform 1 0 16576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_140
timestamp 1698175906
transform 1 0 17024 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_148
timestamp 1698175906
transform 1 0 17920 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_157
timestamp 1698175906
transform 1 0 18928 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698175906
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_123
timestamp 1698175906
transform 1 0 15120 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_153
timestamp 1698175906
transform 1 0 18480 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_169
timestamp 1698175906
transform 1 0 20272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_6
timestamp 1698175906
transform 1 0 2016 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_108
timestamp 1698175906
transform 1 0 13440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita19_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 16576 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18928 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 15568 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 14784 41200 14896 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 41200 16128 42000 16240 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 41200 20160 42000 20272 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 15456 41200 15568 42000 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 19432 27384 19432 27384 0 _000_
rlabel metal2 19992 21336 19992 21336 0 _001_
rlabel metal2 14168 17024 14168 17024 0 _002_
rlabel metal2 21448 14112 21448 14112 0 _003_
rlabel metal2 13944 15456 13944 15456 0 _004_
rlabel metal3 13776 20664 13776 20664 0 _005_
rlabel metal2 24584 21168 24584 21168 0 _006_
rlabel metal2 23688 14840 23688 14840 0 _007_
rlabel metal2 15960 13272 15960 13272 0 _008_
rlabel metal2 15568 28056 15568 28056 0 _009_
rlabel metal3 13664 25704 13664 25704 0 _010_
rlabel metal2 18200 14056 18200 14056 0 _011_
rlabel metal2 21448 25592 21448 25592 0 _012_
rlabel metal2 26264 20328 26264 20328 0 _013_
rlabel metal2 19432 24696 19432 24696 0 _014_
rlabel metal2 16744 14868 16744 14868 0 _015_
rlabel metal2 25424 16184 25424 16184 0 _016_
rlabel metal2 22120 19712 22120 19712 0 _017_
rlabel metal3 13048 20552 13048 20552 0 _018_
rlabel metal3 12992 23016 12992 23016 0 _019_
rlabel metal2 14728 24864 14728 24864 0 _020_
rlabel metal2 23800 25144 23800 25144 0 _021_
rlabel metal2 13160 26656 13160 26656 0 _022_
rlabel metal2 25312 24024 25312 24024 0 _023_
rlabel metal2 25984 17752 25984 17752 0 _024_
rlabel metal2 14728 26936 14728 26936 0 _025_
rlabel metal2 22008 18144 22008 18144 0 _026_
rlabel metal3 20776 18200 20776 18200 0 _027_
rlabel metal2 25984 23912 25984 23912 0 _028_
rlabel metal2 24024 20496 24024 20496 0 _029_
rlabel metal2 27048 17752 27048 17752 0 _030_
rlabel metal2 17976 18144 17976 18144 0 _031_
rlabel metal2 20664 16408 20664 16408 0 _032_
rlabel metal2 19600 20776 19600 20776 0 _033_
rlabel metal2 19096 27720 19096 27720 0 _034_
rlabel metal2 14952 17472 14952 17472 0 _035_
rlabel metal2 18648 18984 18648 18984 0 _036_
rlabel metal2 20104 21224 20104 21224 0 _037_
rlabel metal3 21112 21000 21112 21000 0 _038_
rlabel metal2 14392 18536 14392 18536 0 _039_
rlabel metal2 14728 17696 14728 17696 0 _040_
rlabel metal2 23464 16912 23464 16912 0 _041_
rlabel metal2 22176 14392 22176 14392 0 _042_
rlabel metal2 14504 16464 14504 16464 0 _043_
rlabel metal2 14840 16520 14840 16520 0 _044_
rlabel metal2 14504 20496 14504 20496 0 _045_
rlabel metal3 25816 20664 25816 20664 0 _046_
rlabel metal2 23912 15456 23912 15456 0 _047_
rlabel metal2 18648 14616 18648 14616 0 _048_
rlabel metal2 16856 14280 16856 14280 0 _049_
rlabel metal2 14336 25368 14336 25368 0 _050_
rlabel metal2 15736 27272 15736 27272 0 _051_
rlabel metal2 13720 25088 13720 25088 0 _052_
rlabel metal2 13664 25480 13664 25480 0 _053_
rlabel metal2 19656 13720 19656 13720 0 _054_
rlabel metal2 19320 14448 19320 14448 0 _055_
rlabel metal2 21616 26936 21616 26936 0 _056_
rlabel metal2 23352 19600 23352 19600 0 _057_
rlabel metal2 19432 19040 19432 19040 0 _058_
rlabel metal2 18088 18144 18088 18144 0 _059_
rlabel metal2 14392 23856 14392 23856 0 _060_
rlabel metal2 19040 18536 19040 18536 0 _061_
rlabel metal2 19992 19096 19992 19096 0 _062_
rlabel metal2 17640 22288 17640 22288 0 _063_
rlabel metal3 22512 23912 22512 23912 0 _064_
rlabel metal3 24808 23800 24808 23800 0 _065_
rlabel metal2 25536 19320 25536 19320 0 _066_
rlabel metal2 20776 18760 20776 18760 0 _067_
rlabel metal2 20104 18368 20104 18368 0 _068_
rlabel metal3 19992 23800 19992 23800 0 _069_
rlabel metal3 20776 23688 20776 23688 0 _070_
rlabel metal2 15848 22904 15848 22904 0 _071_
rlabel metal2 21560 21560 21560 21560 0 _072_
rlabel metal2 19880 23912 19880 23912 0 _073_
rlabel metal2 17416 17584 17416 17584 0 _074_
rlabel metal2 18312 19936 18312 19936 0 _075_
rlabel metal2 20328 20608 20328 20608 0 _076_
rlabel metal2 18760 18592 18760 18592 0 _077_
rlabel metal3 18536 15176 18536 15176 0 _078_
rlabel metal2 18872 20384 18872 20384 0 _079_
rlabel metal2 14840 20272 14840 20272 0 _080_
rlabel metal2 23800 21280 23800 21280 0 _081_
rlabel metal2 21224 17248 21224 17248 0 _082_
rlabel metal2 26040 16912 26040 16912 0 _083_
rlabel metal3 16800 20776 16800 20776 0 _084_
rlabel metal2 13832 23576 13832 23576 0 _085_
rlabel metal2 17192 21560 17192 21560 0 _086_
rlabel metal2 14616 22008 14616 22008 0 _087_
rlabel via2 14504 21672 14504 21672 0 _088_
rlabel metal2 13720 24080 13720 24080 0 _089_
rlabel metal2 15288 20440 15288 20440 0 _090_
rlabel metal2 15400 26096 15400 26096 0 _091_
rlabel metal3 21280 22232 21280 22232 0 _092_
rlabel metal2 22792 22680 22792 22680 0 _093_
rlabel metal2 23240 21504 23240 21504 0 _094_
rlabel metal2 23688 24080 23688 24080 0 _095_
rlabel metal2 18256 28504 18256 28504 0 _096_
rlabel metal3 2478 28280 2478 28280 0 clk
rlabel metal2 23464 20776 23464 20776 0 clknet_0_clk
rlabel metal2 22064 14616 22064 14616 0 clknet_1_0__leaf_clk
rlabel metal2 20552 27720 20552 27720 0 clknet_1_1__leaf_clk
rlabel metal2 16352 19320 16352 19320 0 dut19.count\[0\]
rlabel metal3 14616 19208 14616 19208 0 dut19.count\[1\]
rlabel metal2 14952 22736 14952 22736 0 dut19.count\[2\]
rlabel metal2 17024 24584 17024 24584 0 dut19.count\[3\]
rlabel metal2 23576 13552 23576 13552 0 net1
rlabel metal3 18032 28504 18032 28504 0 net10
rlabel metal2 21224 38024 21224 38024 0 net11
rlabel metal2 12040 17192 12040 17192 0 net12
rlabel metal3 12376 20888 12376 20888 0 net13
rlabel metal2 28056 17416 28056 17416 0 net14
rlabel metal2 25256 6356 25256 6356 0 net15
rlabel metal2 17640 5964 17640 5964 0 net16
rlabel metal3 30044 24584 30044 24584 0 net17
rlabel metal2 37912 25928 37912 25928 0 net18
rlabel metal2 27608 16520 27608 16520 0 net19
rlabel metal2 11256 27384 11256 27384 0 net2
rlabel metal2 19096 6356 19096 6356 0 net20
rlabel metal3 33040 19880 33040 19880 0 net21
rlabel metal2 20888 32060 20888 32060 0 net22
rlabel metal3 16184 26936 16184 26936 0 net23
rlabel metal2 15288 29988 15288 29988 0 net24
rlabel metal3 23912 28280 23912 28280 0 net25
rlabel metal3 1246 37016 1246 37016 0 net26
rlabel metal2 21112 5964 21112 5964 0 net3
rlabel metal2 4312 16912 4312 16912 0 net4
rlabel metal3 30380 21672 30380 21672 0 net5
rlabel metal2 37688 25760 37688 25760 0 net6
rlabel metal2 13496 28616 13496 28616 0 net7
rlabel metal2 28168 21504 28168 21504 0 net8
rlabel metal2 25816 25032 25816 25032 0 net9
rlabel metal2 22904 2198 22904 2198 0 segm[10]
rlabel metal3 1358 26936 1358 26936 0 segm[11]
rlabel metal2 20888 2198 20888 2198 0 segm[12]
rlabel metal3 1358 16184 1358 16184 0 segm[13]
rlabel metal2 40040 22344 40040 22344 0 segm[1]
rlabel metal2 39928 25872 39928 25872 0 segm[2]
rlabel metal2 14840 39690 14840 39690 0 segm[3]
rlabel metal2 40040 21504 40040 21504 0 segm[4]
rlabel metal2 40040 23800 40040 23800 0 segm[5]
rlabel metal2 19544 39746 19544 39746 0 segm[6]
rlabel metal2 22232 39746 22232 39746 0 segm[7]
rlabel metal3 1358 16856 1358 16856 0 segm[8]
rlabel metal3 1358 20888 1358 20888 0 segm[9]
rlabel metal3 40642 18200 40642 18200 0 sel[0]
rlabel metal2 24248 2422 24248 2422 0 sel[10]
rlabel metal2 18200 2198 18200 2198 0 sel[11]
rlabel metal2 40040 24360 40040 24360 0 sel[1]
rlabel metal2 40040 25256 40040 25256 0 sel[2]
rlabel metal2 40040 16408 40040 16408 0 sel[3]
rlabel metal2 18872 2422 18872 2422 0 sel[4]
rlabel metal2 40040 20552 40040 20552 0 sel[5]
rlabel metal2 20216 39354 20216 39354 0 sel[6]
rlabel metal2 16184 39354 16184 39354 0 sel[7]
rlabel metal2 15512 38962 15512 38962 0 sel[8]
rlabel metal2 22904 39746 22904 39746 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
