magic
tech gf180mcuD
magscale 1 5
timestamp 1699641753
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 11097 19055 11103 19081
rect 11129 19055 11135 19081
rect 9025 18999 9031 19025
rect 9057 18999 9063 19025
rect 11769 18999 11775 19025
rect 11801 18999 11807 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10375 18745 10401 18751
rect 10375 18713 10401 18719
rect 9865 18607 9871 18633
rect 9897 18607 9903 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 9529 14351 9535 14377
rect 9561 14351 9567 14377
rect 9367 14265 9393 14271
rect 9367 14233 9393 14239
rect 9479 14265 9505 14271
rect 9479 14233 9505 14239
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8689 13903 8695 13929
rect 8721 13903 8727 13929
rect 10649 13903 10655 13929
rect 10681 13903 10687 13929
rect 8471 13873 8497 13879
rect 12391 13873 12417 13879
rect 9081 13847 9087 13873
rect 9113 13847 9119 13873
rect 10145 13847 10151 13873
rect 10177 13847 10183 13873
rect 11041 13847 11047 13873
rect 11073 13847 11079 13873
rect 12105 13847 12111 13873
rect 12137 13847 12143 13873
rect 8471 13841 8497 13847
rect 12391 13841 12417 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 9367 13649 9393 13655
rect 9367 13617 9393 13623
rect 9535 13649 9561 13655
rect 9535 13617 9561 13623
rect 967 13593 993 13599
rect 9759 13593 9785 13599
rect 11663 13593 11689 13599
rect 9193 13567 9199 13593
rect 9225 13567 9231 13593
rect 11097 13567 11103 13593
rect 11129 13567 11135 13593
rect 967 13561 993 13567
rect 9759 13561 9785 13567
rect 11663 13561 11689 13567
rect 11719 13593 11745 13599
rect 11719 13561 11745 13567
rect 10375 13537 10401 13543
rect 11271 13537 11297 13543
rect 2137 13511 2143 13537
rect 2169 13511 2175 13537
rect 7793 13511 7799 13537
rect 7825 13511 7831 13537
rect 10929 13511 10935 13537
rect 10961 13511 10967 13537
rect 10375 13505 10401 13511
rect 11271 13505 11297 13511
rect 7463 13481 7489 13487
rect 9423 13481 9449 13487
rect 10207 13481 10233 13487
rect 8129 13455 8135 13481
rect 8161 13455 8167 13481
rect 10145 13455 10151 13481
rect 10177 13455 10183 13481
rect 7463 13449 7489 13455
rect 9423 13449 9449 13455
rect 10207 13449 10233 13455
rect 10263 13481 10289 13487
rect 10263 13449 10289 13455
rect 11103 13481 11129 13487
rect 11103 13449 11129 13455
rect 11159 13481 11185 13487
rect 11159 13449 11185 13455
rect 11439 13481 11465 13487
rect 11439 13449 11465 13455
rect 11495 13481 11521 13487
rect 11495 13449 11521 13455
rect 7407 13425 7433 13431
rect 7407 13393 7433 13399
rect 10319 13425 10345 13431
rect 10319 13393 10345 13399
rect 20119 13425 20145 13431
rect 20119 13393 20145 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7631 13257 7657 13263
rect 7631 13225 7657 13231
rect 8863 13257 8889 13263
rect 8863 13225 8889 13231
rect 9199 13257 9225 13263
rect 11551 13257 11577 13263
rect 9529 13231 9535 13257
rect 9561 13231 9567 13257
rect 9199 13225 9225 13231
rect 11551 13225 11577 13231
rect 9087 13201 9113 13207
rect 10257 13175 10263 13201
rect 10289 13175 10295 13201
rect 13449 13175 13455 13201
rect 13481 13175 13487 13201
rect 9087 13169 9113 13175
rect 7407 13145 7433 13151
rect 7799 13145 7825 13151
rect 8751 13145 8777 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 6841 13119 6847 13145
rect 6873 13119 6879 13145
rect 7177 13119 7183 13145
rect 7209 13119 7215 13145
rect 7737 13119 7743 13145
rect 7769 13119 7775 13145
rect 7905 13119 7911 13145
rect 7937 13119 7943 13145
rect 7407 13113 7433 13119
rect 7799 13113 7825 13119
rect 8751 13113 8777 13119
rect 8807 13145 8833 13151
rect 8807 13113 8833 13119
rect 9031 13145 9057 13151
rect 9031 13113 9057 13119
rect 9255 13145 9281 13151
rect 9641 13119 9647 13145
rect 9673 13119 9679 13145
rect 9865 13119 9871 13145
rect 9897 13119 9903 13145
rect 12889 13119 12895 13145
rect 12921 13119 12927 13145
rect 13337 13119 13343 13145
rect 13369 13119 13375 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 9255 13113 9281 13119
rect 8135 13089 8161 13095
rect 12783 13089 12809 13095
rect 5777 13063 5783 13089
rect 5809 13063 5815 13089
rect 11321 13063 11327 13089
rect 11353 13063 11359 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 8135 13057 8161 13063
rect 12783 13057 12809 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 7463 13033 7489 13039
rect 7463 13001 7489 13007
rect 12727 13033 12753 13039
rect 12727 13001 12753 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 11327 12865 11353 12871
rect 11327 12833 11353 12839
rect 20007 12809 20033 12815
rect 7345 12783 7351 12809
rect 7377 12783 7383 12809
rect 13449 12783 13455 12809
rect 13481 12783 13487 12809
rect 20007 12777 20033 12783
rect 7407 12753 7433 12759
rect 11489 12727 11495 12753
rect 11521 12727 11527 12753
rect 12049 12727 12055 12753
rect 12081 12727 12087 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 7407 12721 7433 12727
rect 7631 12697 7657 12703
rect 7631 12665 7657 12671
rect 7743 12697 7769 12703
rect 7743 12665 7769 12671
rect 7855 12697 7881 12703
rect 7855 12665 7881 12671
rect 7911 12697 7937 12703
rect 7911 12665 7937 12671
rect 11607 12697 11633 12703
rect 12385 12671 12391 12697
rect 12417 12671 12423 12697
rect 11607 12665 11633 12671
rect 7351 12641 7377 12647
rect 7351 12609 7377 12615
rect 7519 12641 7545 12647
rect 7519 12609 7545 12615
rect 8191 12641 8217 12647
rect 8191 12609 8217 12615
rect 11551 12641 11577 12647
rect 11551 12609 11577 12615
rect 11663 12641 11689 12647
rect 11663 12609 11689 12615
rect 13679 12641 13705 12647
rect 13679 12609 13705 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 6785 12391 6791 12417
rect 6817 12391 6823 12417
rect 9585 12391 9591 12417
rect 9617 12391 9623 12417
rect 12777 12391 12783 12417
rect 12809 12391 12815 12417
rect 9759 12361 9785 12367
rect 7177 12335 7183 12361
rect 7209 12335 7215 12361
rect 9759 12329 9785 12335
rect 10207 12361 10233 12367
rect 10929 12335 10935 12361
rect 10961 12335 10967 12361
rect 12665 12335 12671 12361
rect 12697 12335 12703 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 10207 12329 10233 12335
rect 7407 12305 7433 12311
rect 5721 12279 5727 12305
rect 5753 12279 5759 12305
rect 7407 12273 7433 12279
rect 9983 12305 10009 12311
rect 11265 12279 11271 12305
rect 11297 12279 11303 12305
rect 12329 12279 12335 12305
rect 12361 12279 12367 12305
rect 9983 12273 10009 12279
rect 9927 12249 9953 12255
rect 9927 12217 9953 12223
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 967 12025 993 12031
rect 20007 12025 20033 12031
rect 9921 11999 9927 12025
rect 9953 11999 9959 12025
rect 11377 11999 11383 12025
rect 11409 11999 11415 12025
rect 967 11993 993 11999
rect 20007 11993 20033 11999
rect 10207 11969 10233 11975
rect 11047 11969 11073 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 8465 11943 8471 11969
rect 8497 11943 8503 11969
rect 10761 11943 10767 11969
rect 10793 11943 10799 11969
rect 10207 11937 10233 11943
rect 11047 11937 11073 11943
rect 11159 11969 11185 11975
rect 11159 11937 11185 11943
rect 11271 11969 11297 11975
rect 11887 11969 11913 11975
rect 11713 11943 11719 11969
rect 11745 11943 11751 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 11271 11937 11297 11943
rect 11887 11937 11913 11943
rect 11383 11913 11409 11919
rect 8857 11887 8863 11913
rect 8889 11887 8895 11913
rect 10649 11887 10655 11913
rect 10681 11887 10687 11913
rect 11383 11881 11409 11887
rect 8079 11857 8105 11863
rect 11495 11857 11521 11863
rect 10369 11831 10375 11857
rect 10401 11831 10407 11857
rect 8079 11825 8105 11831
rect 11495 11825 11521 11831
rect 11943 11857 11969 11863
rect 11943 11825 11969 11831
rect 11999 11857 12025 11863
rect 11999 11825 12025 11831
rect 12447 11857 12473 11863
rect 12447 11825 12473 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 8807 11689 8833 11695
rect 8807 11657 8833 11663
rect 10151 11689 10177 11695
rect 10151 11657 10177 11663
rect 14799 11689 14825 11695
rect 14799 11657 14825 11663
rect 8191 11633 8217 11639
rect 7569 11607 7575 11633
rect 7601 11607 7607 11633
rect 8191 11601 8217 11607
rect 8975 11633 9001 11639
rect 9423 11633 9449 11639
rect 9249 11607 9255 11633
rect 9281 11607 9287 11633
rect 10313 11607 10319 11633
rect 10345 11607 10351 11633
rect 10817 11607 10823 11633
rect 10849 11607 10855 11633
rect 8975 11601 9001 11607
rect 9423 11601 9449 11607
rect 8135 11577 8161 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 7905 11551 7911 11577
rect 7937 11551 7943 11577
rect 8135 11545 8161 11551
rect 8247 11577 8273 11583
rect 8247 11545 8273 11551
rect 8415 11577 8441 11583
rect 8415 11545 8441 11551
rect 8751 11577 8777 11583
rect 8751 11545 8777 11551
rect 8863 11577 8889 11583
rect 10655 11577 10681 11583
rect 9809 11551 9815 11577
rect 9841 11551 9847 11577
rect 13113 11551 13119 11577
rect 13145 11551 13151 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 8863 11545 8889 11551
rect 10655 11545 10681 11551
rect 6287 11521 6313 11527
rect 9591 11521 9617 11527
rect 6505 11495 6511 11521
rect 6537 11495 6543 11521
rect 13505 11495 13511 11521
rect 13537 11495 13543 11521
rect 14569 11495 14575 11521
rect 14601 11495 14607 11521
rect 6287 11489 6313 11495
rect 9591 11489 9617 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 6343 11465 6369 11471
rect 6343 11433 6369 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 8191 11297 8217 11303
rect 8191 11265 8217 11271
rect 8695 11241 8721 11247
rect 4937 11215 4943 11241
rect 4969 11215 4975 11241
rect 8695 11209 8721 11215
rect 10599 11241 10625 11247
rect 10599 11209 10625 11215
rect 11383 11241 11409 11247
rect 11383 11209 11409 11215
rect 13455 11241 13481 11247
rect 13455 11209 13481 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 10767 11185 10793 11191
rect 6337 11159 6343 11185
rect 6369 11159 6375 11185
rect 9641 11159 9647 11185
rect 9673 11159 9679 11185
rect 9921 11159 9927 11185
rect 9953 11159 9959 11185
rect 10089 11159 10095 11185
rect 10121 11159 10127 11185
rect 10767 11153 10793 11159
rect 10879 11185 10905 11191
rect 10879 11153 10905 11159
rect 10935 11185 10961 11191
rect 10935 11153 10961 11159
rect 13511 11185 13537 11191
rect 13511 11153 13537 11159
rect 13735 11185 13761 11191
rect 13735 11153 13761 11159
rect 13791 11185 13817 11191
rect 13791 11153 13817 11159
rect 14015 11185 14041 11191
rect 18937 11159 18943 11185
rect 18969 11159 18975 11185
rect 14015 11153 14041 11159
rect 8191 11129 8217 11135
rect 6001 11103 6007 11129
rect 6033 11103 6039 11129
rect 8191 11097 8217 11103
rect 8247 11129 8273 11135
rect 8247 11097 8273 11103
rect 8471 11129 8497 11135
rect 8471 11097 8497 11103
rect 9423 11129 9449 11135
rect 10655 11129 10681 11135
rect 9585 11103 9591 11129
rect 9617 11103 9623 11129
rect 9423 11097 9449 11103
rect 10655 11097 10681 11103
rect 11159 11129 11185 11135
rect 11159 11097 11185 11103
rect 11271 11129 11297 11135
rect 11271 11097 11297 11103
rect 11439 11129 11465 11135
rect 11439 11097 11465 11103
rect 6791 11073 6817 11079
rect 6791 11041 6817 11047
rect 8415 11073 8441 11079
rect 8415 11041 8441 11047
rect 9087 11073 9113 11079
rect 11607 11073 11633 11079
rect 13175 11073 13201 11079
rect 9249 11047 9255 11073
rect 9281 11047 9287 11073
rect 11769 11047 11775 11073
rect 11801 11047 11807 11073
rect 9087 11041 9113 11047
rect 11607 11041 11633 11047
rect 13175 11041 13201 11047
rect 13399 11073 13425 11079
rect 13399 11041 13425 11047
rect 13679 11073 13705 11079
rect 13679 11041 13705 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7351 10905 7377 10911
rect 9025 10879 9031 10905
rect 9057 10879 9063 10905
rect 7351 10873 7377 10879
rect 7183 10849 7209 10855
rect 7183 10817 7209 10823
rect 7799 10849 7825 10855
rect 7799 10817 7825 10823
rect 8079 10849 8105 10855
rect 8079 10817 8105 10823
rect 12671 10849 12697 10855
rect 15297 10823 15303 10849
rect 15329 10823 15335 10849
rect 12671 10817 12697 10823
rect 6959 10793 6985 10799
rect 5329 10767 5335 10793
rect 5361 10767 5367 10793
rect 6959 10761 6985 10767
rect 7015 10793 7041 10799
rect 7407 10793 7433 10799
rect 7289 10767 7295 10793
rect 7321 10767 7327 10793
rect 7015 10761 7041 10767
rect 7407 10761 7433 10767
rect 7575 10793 7601 10799
rect 7575 10761 7601 10767
rect 7911 10793 7937 10799
rect 8863 10793 8889 10799
rect 12615 10793 12641 10799
rect 8185 10767 8191 10793
rect 8217 10767 8223 10793
rect 8297 10767 8303 10793
rect 8329 10767 8335 10793
rect 9193 10767 9199 10793
rect 9225 10767 9231 10793
rect 9529 10767 9535 10793
rect 9561 10767 9567 10793
rect 13561 10767 13567 10793
rect 13593 10767 13599 10793
rect 15185 10767 15191 10793
rect 15217 10767 15223 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 7911 10761 7937 10767
rect 8863 10761 8889 10767
rect 12615 10761 12641 10767
rect 7687 10737 7713 10743
rect 13343 10737 13369 10743
rect 20007 10737 20033 10743
rect 5665 10711 5671 10737
rect 5697 10711 5703 10737
rect 6729 10711 6735 10737
rect 6761 10711 6767 10737
rect 8129 10711 8135 10737
rect 8161 10711 8167 10737
rect 9249 10711 9255 10737
rect 9281 10711 9287 10737
rect 11377 10711 11383 10737
rect 11409 10711 11415 10737
rect 13897 10711 13903 10737
rect 13929 10711 13935 10737
rect 14961 10711 14967 10737
rect 14993 10711 14999 10737
rect 7687 10705 7713 10711
rect 13343 10705 13369 10711
rect 20007 10705 20033 10711
rect 9367 10681 9393 10687
rect 9367 10649 9393 10655
rect 12671 10681 12697 10687
rect 12671 10649 12697 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 6847 10457 6873 10463
rect 20007 10457 20033 10463
rect 7737 10431 7743 10457
rect 7769 10431 7775 10457
rect 13561 10431 13567 10457
rect 13593 10431 13599 10457
rect 6847 10425 6873 10431
rect 20007 10425 20033 10431
rect 7183 10401 7209 10407
rect 10767 10401 10793 10407
rect 14183 10401 14209 10407
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 10985 10375 10991 10401
rect 11017 10375 11023 10401
rect 11377 10375 11383 10401
rect 11409 10375 11415 10401
rect 14905 10375 14911 10401
rect 14937 10375 14943 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 7183 10369 7209 10375
rect 10767 10369 10793 10375
rect 14183 10369 14209 10375
rect 7015 10345 7041 10351
rect 7015 10313 7041 10319
rect 11215 10345 11241 10351
rect 11215 10313 11241 10319
rect 14239 10345 14265 10351
rect 15017 10319 15023 10345
rect 15049 10319 15055 10345
rect 14239 10313 14265 10319
rect 7071 10289 7097 10295
rect 7463 10289 7489 10295
rect 7289 10263 7295 10289
rect 7321 10263 7327 10289
rect 7071 10257 7097 10263
rect 7463 10257 7489 10263
rect 14351 10289 14377 10295
rect 14351 10257 14377 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 13735 10121 13761 10127
rect 7345 10095 7351 10121
rect 7377 10095 7383 10121
rect 8073 10095 8079 10121
rect 8105 10095 8111 10121
rect 8241 10095 8247 10121
rect 8273 10095 8279 10121
rect 10033 10095 10039 10121
rect 10065 10095 10071 10121
rect 13735 10089 13761 10095
rect 7519 10065 7545 10071
rect 12615 10065 12641 10071
rect 9585 10039 9591 10065
rect 9617 10039 9623 10065
rect 9809 10039 9815 10065
rect 9841 10039 9847 10065
rect 10985 10039 10991 10065
rect 11017 10039 11023 10065
rect 11545 10039 11551 10065
rect 11577 10039 11583 10065
rect 7519 10033 7545 10039
rect 12615 10033 12641 10039
rect 13511 10065 13537 10071
rect 13511 10033 13537 10039
rect 13623 10065 13649 10071
rect 13623 10033 13649 10039
rect 12783 10009 12809 10015
rect 7121 9983 7127 10009
rect 7153 9983 7159 10009
rect 7401 9983 7407 10009
rect 7433 9983 7439 10009
rect 7961 9983 7967 10009
rect 7993 9983 7999 10009
rect 8353 9983 8359 10009
rect 8385 9983 8391 10009
rect 9193 9983 9199 10009
rect 9225 9983 9231 10009
rect 9529 9983 9535 10009
rect 9561 9983 9567 10009
rect 10257 9983 10263 10009
rect 10289 9983 10295 10009
rect 11713 9983 11719 10009
rect 11745 9983 11751 10009
rect 12783 9977 12809 9983
rect 12839 10009 12865 10015
rect 12839 9977 12865 9983
rect 13847 10009 13873 10015
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 13847 9977 13873 9983
rect 8975 9953 9001 9959
rect 12671 9953 12697 9959
rect 9137 9927 9143 9953
rect 9169 9927 9175 9953
rect 11321 9927 11327 9953
rect 11353 9927 11359 9953
rect 8975 9921 9001 9927
rect 12671 9921 12697 9927
rect 13343 9953 13369 9959
rect 13343 9921 13369 9927
rect 20007 9953 20033 9959
rect 20007 9921 20033 9927
rect 7233 9871 7239 9897
rect 7265 9871 7271 9897
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8863 9729 8889 9735
rect 8863 9697 8889 9703
rect 967 9673 993 9679
rect 7575 9673 7601 9679
rect 20007 9673 20033 9679
rect 4993 9647 4999 9673
rect 5025 9647 5031 9673
rect 11321 9647 11327 9673
rect 11353 9647 11359 9673
rect 12161 9647 12167 9673
rect 12193 9647 12199 9673
rect 13225 9647 13231 9673
rect 13257 9647 13263 9673
rect 967 9641 993 9647
rect 7575 9641 7601 9647
rect 20007 9641 20033 9647
rect 7239 9617 7265 9623
rect 2137 9591 2143 9617
rect 2169 9591 2175 9617
rect 6449 9591 6455 9617
rect 6481 9591 6487 9617
rect 7177 9591 7183 9617
rect 7209 9591 7215 9617
rect 7239 9585 7265 9591
rect 7631 9617 7657 9623
rect 9087 9617 9113 9623
rect 8409 9591 8415 9617
rect 8441 9591 8447 9617
rect 7631 9585 7657 9591
rect 9087 9585 9113 9591
rect 9983 9617 10009 9623
rect 9983 9585 10009 9591
rect 10151 9617 10177 9623
rect 10151 9585 10177 9591
rect 10655 9617 10681 9623
rect 13735 9617 13761 9623
rect 11489 9591 11495 9617
rect 11521 9591 11527 9617
rect 11825 9591 11831 9617
rect 11857 9591 11863 9617
rect 13393 9591 13399 9617
rect 13425 9591 13431 9617
rect 10655 9585 10681 9591
rect 13735 9585 13761 9591
rect 13847 9617 13873 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 13847 9585 13873 9591
rect 7463 9561 7489 9567
rect 8695 9561 8721 9567
rect 6057 9535 6063 9561
rect 6089 9535 6095 9561
rect 7345 9535 7351 9561
rect 7377 9535 7383 9561
rect 7737 9535 7743 9561
rect 7769 9535 7775 9561
rect 8129 9535 8135 9561
rect 8161 9535 8167 9561
rect 8521 9535 8527 9561
rect 8553 9535 8559 9561
rect 7463 9529 7489 9535
rect 8695 9529 8721 9535
rect 8919 9561 8945 9567
rect 13567 9561 13593 9567
rect 9249 9535 9255 9561
rect 9281 9535 9287 9561
rect 10817 9535 10823 9561
rect 10849 9535 10855 9561
rect 8919 9529 8945 9535
rect 13567 9529 13593 9535
rect 14239 9561 14265 9567
rect 14239 9529 14265 9535
rect 6791 9505 6817 9511
rect 8807 9505 8833 9511
rect 7233 9479 7239 9505
rect 7265 9479 7271 9505
rect 6791 9473 6817 9479
rect 8807 9473 8833 9479
rect 10039 9505 10065 9511
rect 10039 9473 10065 9479
rect 13511 9505 13537 9511
rect 13511 9473 13537 9479
rect 13791 9505 13817 9511
rect 13791 9473 13817 9479
rect 13959 9505 13985 9511
rect 13959 9473 13985 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 7127 9337 7153 9343
rect 10991 9337 11017 9343
rect 10761 9311 10767 9337
rect 10793 9311 10799 9337
rect 7127 9305 7153 9311
rect 10991 9305 11017 9311
rect 13007 9337 13033 9343
rect 13007 9305 13033 9311
rect 7519 9281 7545 9287
rect 10935 9281 10961 9287
rect 7401 9255 7407 9281
rect 7433 9255 7439 9281
rect 10201 9255 10207 9281
rect 10233 9255 10239 9281
rect 11881 9255 11887 9281
rect 11913 9255 11919 9281
rect 13617 9255 13623 9281
rect 13649 9255 13655 9281
rect 7519 9249 7545 9255
rect 10935 9249 10961 9255
rect 6735 9225 6761 9231
rect 6735 9193 6761 9199
rect 6959 9225 6985 9231
rect 7295 9225 7321 9231
rect 8695 9225 8721 9231
rect 7233 9199 7239 9225
rect 7265 9199 7271 9225
rect 8129 9199 8135 9225
rect 8161 9199 8167 9225
rect 6959 9193 6985 9199
rect 7295 9193 7321 9199
rect 8695 9193 8721 9199
rect 8975 9225 9001 9231
rect 10599 9225 10625 9231
rect 10089 9199 10095 9225
rect 10121 9199 10127 9225
rect 8975 9193 9001 9199
rect 10599 9193 10625 9199
rect 11719 9225 11745 9231
rect 11719 9193 11745 9199
rect 12951 9225 12977 9231
rect 13281 9199 13287 9225
rect 13313 9199 13319 9225
rect 12951 9193 12977 9199
rect 6679 9169 6705 9175
rect 6679 9137 6705 9143
rect 6903 9169 6929 9175
rect 6903 9137 6929 9143
rect 7855 9169 7881 9175
rect 12335 9169 12361 9175
rect 8185 9143 8191 9169
rect 8217 9143 8223 9169
rect 14681 9143 14687 9169
rect 14713 9143 14719 9169
rect 7855 9137 7881 9143
rect 12335 9137 12361 9143
rect 10991 9113 11017 9119
rect 10991 9081 11017 9087
rect 12839 9113 12865 9119
rect 12839 9081 12865 9087
rect 13007 9113 13033 9119
rect 13007 9081 13033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 8247 8945 8273 8951
rect 11887 8945 11913 8951
rect 8409 8919 8415 8945
rect 8441 8919 8447 8945
rect 8247 8913 8273 8919
rect 11887 8913 11913 8919
rect 8135 8889 8161 8895
rect 20007 8889 20033 8895
rect 7345 8863 7351 8889
rect 7377 8863 7383 8889
rect 13225 8863 13231 8889
rect 13257 8863 13263 8889
rect 14289 8863 14295 8889
rect 14321 8863 14327 8889
rect 8135 8857 8161 8863
rect 20007 8857 20033 8863
rect 7743 8833 7769 8839
rect 7065 8807 7071 8833
rect 7097 8807 7103 8833
rect 7743 8801 7769 8807
rect 8583 8833 8609 8839
rect 8583 8801 8609 8807
rect 10823 8833 10849 8839
rect 14631 8833 14657 8839
rect 11881 8807 11887 8833
rect 11913 8807 11919 8833
rect 12889 8807 12895 8833
rect 12921 8807 12927 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 10823 8801 10849 8807
rect 14631 8801 14657 8807
rect 11719 8777 11745 8783
rect 7905 8751 7911 8777
rect 7937 8751 7943 8777
rect 8745 8751 8751 8777
rect 8777 8751 8783 8777
rect 11719 8745 11745 8751
rect 6959 8721 6985 8727
rect 6959 8689 6985 8695
rect 7575 8721 7601 8727
rect 10649 8695 10655 8721
rect 10681 8695 10687 8721
rect 7575 8689 7601 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 8247 8553 8273 8559
rect 7233 8527 7239 8553
rect 7265 8527 7271 8553
rect 7905 8527 7911 8553
rect 7937 8527 7943 8553
rect 8247 8521 8273 8527
rect 9311 8553 9337 8559
rect 9311 8521 9337 8527
rect 9423 8553 9449 8559
rect 9423 8521 9449 8527
rect 10711 8553 10737 8559
rect 10711 8521 10737 8527
rect 11551 8553 11577 8559
rect 11551 8521 11577 8527
rect 11607 8553 11633 8559
rect 11607 8521 11633 8527
rect 7631 8497 7657 8503
rect 5833 8471 5839 8497
rect 5865 8471 5871 8497
rect 7631 8465 7657 8471
rect 9815 8497 9841 8503
rect 9815 8465 9841 8471
rect 9927 8497 9953 8503
rect 9927 8465 9953 8471
rect 11103 8497 11129 8503
rect 11663 8497 11689 8503
rect 11209 8471 11215 8497
rect 11241 8471 11247 8497
rect 11103 8465 11129 8471
rect 11663 8465 11689 8471
rect 13399 8497 13425 8503
rect 13399 8465 13425 8471
rect 8079 8441 8105 8447
rect 5497 8415 5503 8441
rect 5529 8415 5535 8441
rect 7345 8415 7351 8441
rect 7377 8415 7383 8441
rect 8079 8409 8105 8415
rect 9591 8441 9617 8447
rect 9591 8409 9617 8415
rect 10151 8441 10177 8447
rect 10599 8441 10625 8447
rect 10425 8415 10431 8441
rect 10457 8415 10463 8441
rect 10151 8409 10177 8415
rect 10599 8409 10625 8415
rect 10879 8441 10905 8447
rect 10879 8409 10905 8415
rect 11271 8441 11297 8447
rect 11271 8409 11297 8415
rect 11327 8441 11353 8447
rect 11769 8415 11775 8441
rect 11801 8415 11807 8441
rect 11881 8415 11887 8441
rect 11913 8415 11919 8441
rect 13561 8415 13567 8441
rect 13593 8415 13599 8441
rect 11327 8409 11353 8415
rect 10039 8385 10065 8391
rect 6897 8359 6903 8385
rect 6929 8359 6935 8385
rect 10039 8353 10065 8359
rect 10655 8385 10681 8391
rect 10655 8353 10681 8359
rect 10935 8385 10961 8391
rect 10935 8353 10961 8359
rect 13455 8385 13481 8391
rect 13455 8353 13481 8359
rect 7743 8329 7769 8335
rect 7743 8297 7769 8303
rect 9255 8329 9281 8335
rect 9255 8297 9281 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 7743 8161 7769 8167
rect 7743 8129 7769 8135
rect 9311 8161 9337 8167
rect 9311 8129 9337 8135
rect 9423 8161 9449 8167
rect 9423 8129 9449 8135
rect 9535 8161 9561 8167
rect 9535 8129 9561 8135
rect 9815 8161 9841 8167
rect 9815 8129 9841 8135
rect 9927 8161 9953 8167
rect 9927 8129 9953 8135
rect 11719 8161 11745 8167
rect 11719 8129 11745 8135
rect 11775 8161 11801 8167
rect 11775 8129 11801 8135
rect 10039 8105 10065 8111
rect 9081 8079 9087 8105
rect 9113 8079 9119 8105
rect 10039 8073 10065 8079
rect 8695 8049 8721 8055
rect 9591 8049 9617 8055
rect 9025 8023 9031 8049
rect 9057 8023 9063 8049
rect 8695 8017 8721 8023
rect 9591 8017 9617 8023
rect 10151 8049 10177 8055
rect 10151 8017 10177 8023
rect 11607 8049 11633 8055
rect 11607 8017 11633 8023
rect 12559 8049 12585 8055
rect 12559 8017 12585 8023
rect 7631 7993 7657 7999
rect 7631 7961 7657 7967
rect 8807 7993 8833 7999
rect 8807 7961 8833 7967
rect 8863 7993 8889 7999
rect 8863 7961 8889 7967
rect 11999 7993 12025 7999
rect 11999 7961 12025 7967
rect 12111 7993 12137 7999
rect 12111 7961 12137 7967
rect 12279 7993 12305 7999
rect 12279 7961 12305 7967
rect 12391 7993 12417 7999
rect 12391 7961 12417 7967
rect 7015 7937 7041 7943
rect 7015 7905 7041 7911
rect 7687 7937 7713 7943
rect 7687 7905 7713 7911
rect 9367 7937 9393 7943
rect 9367 7905 9393 7911
rect 10207 7937 10233 7943
rect 10207 7905 10233 7911
rect 10263 7937 10289 7943
rect 10263 7905 10289 7911
rect 11775 7937 11801 7943
rect 11775 7905 11801 7911
rect 12167 7937 12193 7943
rect 12167 7905 12193 7911
rect 12503 7937 12529 7943
rect 12503 7905 12529 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 9087 7713 9113 7719
rect 6673 7687 6679 7713
rect 6705 7687 6711 7713
rect 9087 7681 9113 7687
rect 9143 7713 9169 7719
rect 9143 7681 9169 7687
rect 9255 7713 9281 7719
rect 9255 7681 9281 7687
rect 9367 7713 9393 7719
rect 9367 7681 9393 7687
rect 10319 7713 10345 7719
rect 10319 7681 10345 7687
rect 10375 7713 10401 7719
rect 11265 7687 11271 7713
rect 11297 7687 11303 7713
rect 10375 7681 10401 7687
rect 10095 7657 10121 7663
rect 6337 7631 6343 7657
rect 6369 7631 6375 7657
rect 10095 7625 10121 7631
rect 10207 7657 10233 7663
rect 12671 7657 12697 7663
rect 10929 7631 10935 7657
rect 10961 7631 10967 7657
rect 10207 7625 10233 7631
rect 12671 7625 12697 7631
rect 7967 7601 7993 7607
rect 7737 7575 7743 7601
rect 7769 7575 7775 7601
rect 7967 7569 7993 7575
rect 8751 7601 8777 7607
rect 12329 7575 12335 7601
rect 12361 7575 12367 7601
rect 8751 7569 8777 7575
rect 10487 7545 10513 7551
rect 10487 7513 10513 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 13287 7321 13313 7327
rect 7681 7295 7687 7321
rect 7713 7295 7719 7321
rect 8745 7295 8751 7321
rect 8777 7295 8783 7321
rect 9305 7295 9311 7321
rect 9337 7295 9343 7321
rect 10369 7295 10375 7321
rect 10401 7295 10407 7321
rect 11937 7295 11943 7321
rect 11969 7295 11975 7321
rect 13001 7295 13007 7321
rect 13033 7295 13039 7321
rect 13287 7289 13313 7295
rect 7345 7239 7351 7265
rect 7377 7239 7383 7265
rect 8913 7239 8919 7265
rect 8945 7239 8951 7265
rect 11545 7239 11551 7265
rect 11577 7239 11583 7265
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8919 6985 8945 6991
rect 8919 6953 8945 6959
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9529 2143 9535 2169
rect 9561 2143 9567 2169
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 10039 2057 10065 2063
rect 10039 2025 10065 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 11047 1833 11073 1839
rect 11047 1801 11073 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 10537 1751 10543 1777
rect 10569 1751 10575 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 10095 1665 10121 1671
rect 10095 1633 10121 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 12783 19111 12809 19137
rect 11103 19055 11129 19081
rect 9031 18999 9057 19025
rect 11775 18999 11801 19025
rect 12279 18999 12305 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10375 18719 10401 18745
rect 9871 18607 9897 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9535 14351 9561 14377
rect 9367 14239 9393 14265
rect 9479 14239 9505 14265
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8695 13903 8721 13929
rect 10655 13903 10681 13929
rect 8471 13847 8497 13873
rect 9087 13847 9113 13873
rect 10151 13847 10177 13873
rect 11047 13847 11073 13873
rect 12111 13847 12137 13873
rect 12391 13847 12417 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9367 13623 9393 13649
rect 9535 13623 9561 13649
rect 967 13567 993 13593
rect 9199 13567 9225 13593
rect 9759 13567 9785 13593
rect 11103 13567 11129 13593
rect 11663 13567 11689 13593
rect 11719 13567 11745 13593
rect 2143 13511 2169 13537
rect 7799 13511 7825 13537
rect 10375 13511 10401 13537
rect 10935 13511 10961 13537
rect 11271 13511 11297 13537
rect 7463 13455 7489 13481
rect 8135 13455 8161 13481
rect 9423 13455 9449 13481
rect 10151 13455 10177 13481
rect 10207 13455 10233 13481
rect 10263 13455 10289 13481
rect 11103 13455 11129 13481
rect 11159 13455 11185 13481
rect 11439 13455 11465 13481
rect 11495 13455 11521 13481
rect 7407 13399 7433 13425
rect 10319 13399 10345 13425
rect 20119 13399 20145 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7631 13231 7657 13257
rect 8863 13231 8889 13257
rect 9199 13231 9225 13257
rect 9535 13231 9561 13257
rect 11551 13231 11577 13257
rect 9087 13175 9113 13201
rect 10263 13175 10289 13201
rect 13455 13175 13481 13201
rect 2143 13119 2169 13145
rect 6847 13119 6873 13145
rect 7183 13119 7209 13145
rect 7407 13119 7433 13145
rect 7743 13119 7769 13145
rect 7799 13119 7825 13145
rect 7911 13119 7937 13145
rect 8751 13119 8777 13145
rect 8807 13119 8833 13145
rect 9031 13119 9057 13145
rect 9255 13119 9281 13145
rect 9647 13119 9673 13145
rect 9871 13119 9897 13145
rect 12895 13119 12921 13145
rect 13343 13119 13369 13145
rect 18831 13119 18857 13145
rect 5783 13063 5809 13089
rect 8135 13063 8161 13089
rect 11327 13063 11353 13089
rect 12783 13063 12809 13089
rect 19951 13063 19977 13089
rect 967 13007 993 13033
rect 7463 13007 7489 13033
rect 12727 13007 12753 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 11327 12839 11353 12865
rect 7351 12783 7377 12809
rect 13455 12783 13481 12809
rect 20007 12783 20033 12809
rect 7407 12727 7433 12753
rect 11495 12727 11521 12753
rect 12055 12727 12081 12753
rect 18831 12727 18857 12753
rect 7631 12671 7657 12697
rect 7743 12671 7769 12697
rect 7855 12671 7881 12697
rect 7911 12671 7937 12697
rect 11607 12671 11633 12697
rect 12391 12671 12417 12697
rect 7351 12615 7377 12641
rect 7519 12615 7545 12641
rect 8191 12615 8217 12641
rect 11551 12615 11577 12641
rect 11663 12615 11689 12641
rect 13679 12615 13705 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 6791 12391 6817 12417
rect 9591 12391 9617 12417
rect 12783 12391 12809 12417
rect 7183 12335 7209 12361
rect 9759 12335 9785 12361
rect 10207 12335 10233 12361
rect 10935 12335 10961 12361
rect 12671 12335 12697 12361
rect 18831 12335 18857 12361
rect 5727 12279 5753 12305
rect 7407 12279 7433 12305
rect 9983 12279 10009 12305
rect 11271 12279 11297 12305
rect 12335 12279 12361 12305
rect 9927 12223 9953 12249
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 967 11999 993 12025
rect 9927 11999 9953 12025
rect 11383 11999 11409 12025
rect 20007 11999 20033 12025
rect 2143 11943 2169 11969
rect 8471 11943 8497 11969
rect 10207 11943 10233 11969
rect 10767 11943 10793 11969
rect 11047 11943 11073 11969
rect 11159 11943 11185 11969
rect 11271 11943 11297 11969
rect 11719 11943 11745 11969
rect 11887 11943 11913 11969
rect 18831 11943 18857 11969
rect 8863 11887 8889 11913
rect 10655 11887 10681 11913
rect 11383 11887 11409 11913
rect 8079 11831 8105 11857
rect 10375 11831 10401 11857
rect 11495 11831 11521 11857
rect 11943 11831 11969 11857
rect 11999 11831 12025 11857
rect 12447 11831 12473 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 8807 11663 8833 11689
rect 10151 11663 10177 11689
rect 14799 11663 14825 11689
rect 7575 11607 7601 11633
rect 8191 11607 8217 11633
rect 8975 11607 9001 11633
rect 9255 11607 9281 11633
rect 9423 11607 9449 11633
rect 10319 11607 10345 11633
rect 10823 11607 10849 11633
rect 2143 11551 2169 11577
rect 7911 11551 7937 11577
rect 8135 11551 8161 11577
rect 8247 11551 8273 11577
rect 8415 11551 8441 11577
rect 8751 11551 8777 11577
rect 8863 11551 8889 11577
rect 9815 11551 9841 11577
rect 10655 11551 10681 11577
rect 13119 11551 13145 11577
rect 18831 11551 18857 11577
rect 6287 11495 6313 11521
rect 6511 11495 6537 11521
rect 9591 11495 9617 11521
rect 13511 11495 13537 11521
rect 14575 11495 14601 11521
rect 967 11439 993 11465
rect 6343 11439 6369 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 8191 11271 8217 11297
rect 4943 11215 4969 11241
rect 8695 11215 8721 11241
rect 10599 11215 10625 11241
rect 11383 11215 11409 11241
rect 13455 11215 13481 11241
rect 20007 11215 20033 11241
rect 6343 11159 6369 11185
rect 9647 11159 9673 11185
rect 9927 11159 9953 11185
rect 10095 11159 10121 11185
rect 10767 11159 10793 11185
rect 10879 11159 10905 11185
rect 10935 11159 10961 11185
rect 13511 11159 13537 11185
rect 13735 11159 13761 11185
rect 13791 11159 13817 11185
rect 14015 11159 14041 11185
rect 18943 11159 18969 11185
rect 6007 11103 6033 11129
rect 8191 11103 8217 11129
rect 8247 11103 8273 11129
rect 8471 11103 8497 11129
rect 9423 11103 9449 11129
rect 9591 11103 9617 11129
rect 10655 11103 10681 11129
rect 11159 11103 11185 11129
rect 11271 11103 11297 11129
rect 11439 11103 11465 11129
rect 6791 11047 6817 11073
rect 8415 11047 8441 11073
rect 9087 11047 9113 11073
rect 9255 11047 9281 11073
rect 11607 11047 11633 11073
rect 11775 11047 11801 11073
rect 13175 11047 13201 11073
rect 13399 11047 13425 11073
rect 13679 11047 13705 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7351 10879 7377 10905
rect 9031 10879 9057 10905
rect 7183 10823 7209 10849
rect 7799 10823 7825 10849
rect 8079 10823 8105 10849
rect 12671 10823 12697 10849
rect 15303 10823 15329 10849
rect 5335 10767 5361 10793
rect 6959 10767 6985 10793
rect 7015 10767 7041 10793
rect 7295 10767 7321 10793
rect 7407 10767 7433 10793
rect 7575 10767 7601 10793
rect 7911 10767 7937 10793
rect 8191 10767 8217 10793
rect 8303 10767 8329 10793
rect 8863 10767 8889 10793
rect 9199 10767 9225 10793
rect 9535 10767 9561 10793
rect 12615 10767 12641 10793
rect 13567 10767 13593 10793
rect 15191 10767 15217 10793
rect 18831 10767 18857 10793
rect 5671 10711 5697 10737
rect 6735 10711 6761 10737
rect 7687 10711 7713 10737
rect 8135 10711 8161 10737
rect 9255 10711 9281 10737
rect 11383 10711 11409 10737
rect 13343 10711 13369 10737
rect 13903 10711 13929 10737
rect 14967 10711 14993 10737
rect 20007 10711 20033 10737
rect 9367 10655 9393 10681
rect 12671 10655 12697 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 6847 10431 6873 10457
rect 7743 10431 7769 10457
rect 13567 10431 13593 10457
rect 20007 10431 20033 10457
rect 7183 10375 7209 10401
rect 10039 10375 10065 10401
rect 10767 10375 10793 10401
rect 10991 10375 11017 10401
rect 11383 10375 11409 10401
rect 14183 10375 14209 10401
rect 14911 10375 14937 10401
rect 18831 10375 18857 10401
rect 7015 10319 7041 10345
rect 11215 10319 11241 10345
rect 14239 10319 14265 10345
rect 15023 10319 15049 10345
rect 7071 10263 7097 10289
rect 7295 10263 7321 10289
rect 7463 10263 7489 10289
rect 14351 10263 14377 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7351 10095 7377 10121
rect 8079 10095 8105 10121
rect 8247 10095 8273 10121
rect 10039 10095 10065 10121
rect 13735 10095 13761 10121
rect 7519 10039 7545 10065
rect 9591 10039 9617 10065
rect 9815 10039 9841 10065
rect 10991 10039 11017 10065
rect 11551 10039 11577 10065
rect 12615 10039 12641 10065
rect 13511 10039 13537 10065
rect 13623 10039 13649 10065
rect 7127 9983 7153 10009
rect 7407 9983 7433 10009
rect 7967 9983 7993 10009
rect 8359 9983 8385 10009
rect 9199 9983 9225 10009
rect 9535 9983 9561 10009
rect 10263 9983 10289 10009
rect 11719 9983 11745 10009
rect 12783 9983 12809 10009
rect 12839 9983 12865 10009
rect 13847 9983 13873 10009
rect 18831 9983 18857 10009
rect 8975 9927 9001 9953
rect 9143 9927 9169 9953
rect 11327 9927 11353 9953
rect 12671 9927 12697 9953
rect 13343 9927 13369 9953
rect 20007 9927 20033 9953
rect 7239 9871 7265 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8863 9703 8889 9729
rect 967 9647 993 9673
rect 4999 9647 5025 9673
rect 7575 9647 7601 9673
rect 11327 9647 11353 9673
rect 12167 9647 12193 9673
rect 13231 9647 13257 9673
rect 20007 9647 20033 9673
rect 2143 9591 2169 9617
rect 6455 9591 6481 9617
rect 7183 9591 7209 9617
rect 7239 9591 7265 9617
rect 7631 9591 7657 9617
rect 8415 9591 8441 9617
rect 9087 9591 9113 9617
rect 9983 9591 10009 9617
rect 10151 9591 10177 9617
rect 10655 9591 10681 9617
rect 11495 9591 11521 9617
rect 11831 9591 11857 9617
rect 13399 9591 13425 9617
rect 13735 9591 13761 9617
rect 13847 9591 13873 9617
rect 18831 9591 18857 9617
rect 6063 9535 6089 9561
rect 7351 9535 7377 9561
rect 7463 9535 7489 9561
rect 7743 9535 7769 9561
rect 8135 9535 8161 9561
rect 8527 9535 8553 9561
rect 8695 9535 8721 9561
rect 8919 9535 8945 9561
rect 9255 9535 9281 9561
rect 10823 9535 10849 9561
rect 13567 9535 13593 9561
rect 14239 9535 14265 9561
rect 6791 9479 6817 9505
rect 7239 9479 7265 9505
rect 8807 9479 8833 9505
rect 10039 9479 10065 9505
rect 13511 9479 13537 9505
rect 13791 9479 13817 9505
rect 13959 9479 13985 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7127 9311 7153 9337
rect 10767 9311 10793 9337
rect 10991 9311 11017 9337
rect 13007 9311 13033 9337
rect 7407 9255 7433 9281
rect 7519 9255 7545 9281
rect 10207 9255 10233 9281
rect 10935 9255 10961 9281
rect 11887 9255 11913 9281
rect 13623 9255 13649 9281
rect 6735 9199 6761 9225
rect 6959 9199 6985 9225
rect 7239 9199 7265 9225
rect 7295 9199 7321 9225
rect 8135 9199 8161 9225
rect 8695 9199 8721 9225
rect 8975 9199 9001 9225
rect 10095 9199 10121 9225
rect 10599 9199 10625 9225
rect 11719 9199 11745 9225
rect 12951 9199 12977 9225
rect 13287 9199 13313 9225
rect 6679 9143 6705 9169
rect 6903 9143 6929 9169
rect 7855 9143 7881 9169
rect 8191 9143 8217 9169
rect 12335 9143 12361 9169
rect 14687 9143 14713 9169
rect 10991 9087 11017 9113
rect 12839 9087 12865 9113
rect 13007 9087 13033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 8247 8919 8273 8945
rect 8415 8919 8441 8945
rect 11887 8919 11913 8945
rect 7351 8863 7377 8889
rect 8135 8863 8161 8889
rect 13231 8863 13257 8889
rect 14295 8863 14321 8889
rect 20007 8863 20033 8889
rect 7071 8807 7097 8833
rect 7743 8807 7769 8833
rect 8583 8807 8609 8833
rect 10823 8807 10849 8833
rect 11887 8807 11913 8833
rect 12895 8807 12921 8833
rect 14631 8807 14657 8833
rect 18831 8807 18857 8833
rect 7911 8751 7937 8777
rect 8751 8751 8777 8777
rect 11719 8751 11745 8777
rect 6959 8695 6985 8721
rect 7575 8695 7601 8721
rect 10655 8695 10681 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7239 8527 7265 8553
rect 7911 8527 7937 8553
rect 8247 8527 8273 8553
rect 9311 8527 9337 8553
rect 9423 8527 9449 8553
rect 10711 8527 10737 8553
rect 11551 8527 11577 8553
rect 11607 8527 11633 8553
rect 5839 8471 5865 8497
rect 7631 8471 7657 8497
rect 9815 8471 9841 8497
rect 9927 8471 9953 8497
rect 11103 8471 11129 8497
rect 11215 8471 11241 8497
rect 11663 8471 11689 8497
rect 13399 8471 13425 8497
rect 5503 8415 5529 8441
rect 7351 8415 7377 8441
rect 8079 8415 8105 8441
rect 9591 8415 9617 8441
rect 10151 8415 10177 8441
rect 10431 8415 10457 8441
rect 10599 8415 10625 8441
rect 10879 8415 10905 8441
rect 11271 8415 11297 8441
rect 11327 8415 11353 8441
rect 11775 8415 11801 8441
rect 11887 8415 11913 8441
rect 13567 8415 13593 8441
rect 6903 8359 6929 8385
rect 10039 8359 10065 8385
rect 10655 8359 10681 8385
rect 10935 8359 10961 8385
rect 13455 8359 13481 8385
rect 7743 8303 7769 8329
rect 9255 8303 9281 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 7743 8135 7769 8161
rect 9311 8135 9337 8161
rect 9423 8135 9449 8161
rect 9535 8135 9561 8161
rect 9815 8135 9841 8161
rect 9927 8135 9953 8161
rect 11719 8135 11745 8161
rect 11775 8135 11801 8161
rect 9087 8079 9113 8105
rect 10039 8079 10065 8105
rect 8695 8023 8721 8049
rect 9031 8023 9057 8049
rect 9591 8023 9617 8049
rect 10151 8023 10177 8049
rect 11607 8023 11633 8049
rect 12559 8023 12585 8049
rect 7631 7967 7657 7993
rect 8807 7967 8833 7993
rect 8863 7967 8889 7993
rect 11999 7967 12025 7993
rect 12111 7967 12137 7993
rect 12279 7967 12305 7993
rect 12391 7967 12417 7993
rect 7015 7911 7041 7937
rect 7687 7911 7713 7937
rect 9367 7911 9393 7937
rect 10207 7911 10233 7937
rect 10263 7911 10289 7937
rect 11775 7911 11801 7937
rect 12167 7911 12193 7937
rect 12503 7911 12529 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 6679 7687 6705 7713
rect 9087 7687 9113 7713
rect 9143 7687 9169 7713
rect 9255 7687 9281 7713
rect 9367 7687 9393 7713
rect 10319 7687 10345 7713
rect 10375 7687 10401 7713
rect 11271 7687 11297 7713
rect 6343 7631 6369 7657
rect 10095 7631 10121 7657
rect 10207 7631 10233 7657
rect 10935 7631 10961 7657
rect 12671 7631 12697 7657
rect 7743 7575 7769 7601
rect 7967 7575 7993 7601
rect 8751 7575 8777 7601
rect 12335 7575 12361 7601
rect 10487 7519 10513 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 7687 7295 7713 7321
rect 8751 7295 8777 7321
rect 9311 7295 9337 7321
rect 10375 7295 10401 7321
rect 11943 7295 11969 7321
rect 13007 7295 13033 7321
rect 13287 7295 13313 7321
rect 7351 7239 7377 7265
rect 8919 7239 8945 7265
rect 11551 7239 11577 7265
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8919 6959 8945 6985
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9535 2143 9561 2169
rect 12615 2143 12641 2169
rect 10039 2031 10065 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 11047 1807 11073 1833
rect 12783 1807 12809 1833
rect 10543 1751 10569 1777
rect 12279 1751 12305 1777
rect 10095 1639 10121 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 9072 20600 9128 21000
rect 9744 20600 9800 21000
rect 11088 20600 11144 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 9086 19138 9114 20600
rect 9310 19138 9338 19143
rect 9086 19137 9338 19138
rect 9086 19111 9311 19137
rect 9337 19111 9338 19137
rect 9086 19110 9338 19111
rect 9310 19105 9338 19110
rect 9030 19025 9058 19031
rect 9030 18999 9031 19025
rect 9057 18999 9058 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 8750 14266 8778 14271
rect 8694 13929 8722 13935
rect 8694 13903 8695 13929
rect 8721 13903 8722 13929
rect 8470 13874 8498 13879
rect 8694 13874 8722 13903
rect 8358 13873 8722 13874
rect 8358 13847 8471 13873
rect 8497 13847 8722 13873
rect 8358 13846 8722 13847
rect 2086 13818 2114 13823
rect 966 13593 994 13599
rect 966 13567 967 13593
rect 993 13567 994 13593
rect 966 13146 994 13567
rect 966 13113 994 13118
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 2086 11074 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 2142 13537 2170 13543
rect 2142 13511 2143 13537
rect 2169 13511 2170 13537
rect 2142 13482 2170 13511
rect 7798 13537 7826 13543
rect 7798 13511 7799 13537
rect 7825 13511 7826 13537
rect 2142 13449 2170 13454
rect 5782 13482 5810 13487
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 5726 13146 5754 13151
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 5726 12698 5754 13118
rect 5782 13089 5810 13454
rect 7462 13482 7490 13487
rect 7462 13435 7490 13454
rect 7798 13454 7826 13511
rect 8134 13481 8162 13487
rect 8134 13455 8135 13481
rect 8161 13455 8162 13481
rect 7406 13425 7434 13431
rect 7406 13399 7407 13425
rect 7433 13399 7434 13425
rect 6846 13146 6874 13151
rect 6846 13099 6874 13118
rect 7182 13145 7210 13151
rect 7182 13119 7183 13145
rect 7209 13119 7210 13145
rect 5782 13063 5783 13089
rect 5809 13063 5810 13089
rect 5782 13057 5810 13063
rect 6902 12754 6930 12759
rect 5726 12305 5754 12670
rect 6790 12726 6902 12754
rect 6790 12417 6818 12726
rect 6902 12721 6930 12726
rect 6790 12391 6791 12417
rect 6817 12391 6818 12417
rect 6790 12385 6818 12391
rect 5726 12279 5727 12305
rect 5753 12279 5754 12305
rect 5726 12273 5754 12279
rect 7182 12361 7210 13119
rect 7406 13145 7434 13399
rect 7630 13426 7658 13431
rect 7798 13426 8106 13454
rect 7630 13257 7658 13398
rect 7630 13231 7631 13257
rect 7657 13231 7658 13257
rect 7630 13225 7658 13231
rect 7406 13119 7407 13145
rect 7433 13119 7434 13145
rect 7406 13113 7434 13119
rect 7742 13145 7770 13151
rect 7742 13119 7743 13145
rect 7769 13119 7770 13145
rect 7742 13090 7770 13119
rect 7798 13146 7826 13151
rect 7798 13099 7826 13118
rect 7910 13145 7938 13151
rect 7910 13119 7911 13145
rect 7937 13119 7938 13145
rect 7462 13034 7490 13039
rect 7350 12809 7378 12815
rect 7350 12783 7351 12809
rect 7377 12783 7378 12809
rect 7350 12754 7378 12783
rect 7350 12721 7378 12726
rect 7406 12810 7434 12815
rect 7406 12753 7434 12782
rect 7406 12727 7407 12753
rect 7433 12727 7434 12753
rect 7406 12721 7434 12727
rect 7350 12642 7378 12647
rect 7350 12595 7378 12614
rect 7182 12335 7183 12361
rect 7209 12335 7210 12361
rect 7182 12306 7210 12335
rect 7406 12306 7434 12311
rect 7182 12305 7434 12306
rect 7182 12279 7407 12305
rect 7433 12279 7434 12305
rect 7182 12278 7434 12279
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 6510 11970 6538 11975
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 4942 11522 4970 11527
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 4942 11241 4970 11494
rect 6286 11522 6314 11527
rect 6286 11475 6314 11494
rect 6510 11521 6538 11942
rect 6510 11495 6511 11521
rect 6537 11495 6538 11521
rect 6342 11466 6370 11471
rect 6342 11465 6426 11466
rect 6342 11439 6343 11465
rect 6369 11439 6426 11465
rect 6342 11438 6426 11439
rect 6342 11433 6370 11438
rect 4942 11215 4943 11241
rect 4969 11215 4970 11241
rect 4942 11209 4970 11215
rect 6342 11185 6370 11191
rect 6342 11159 6343 11185
rect 6369 11159 6370 11185
rect 2086 11041 2114 11046
rect 6006 11129 6034 11135
rect 6006 11103 6007 11129
rect 6033 11103 6034 11129
rect 5334 10906 5362 10911
rect 5334 10793 5362 10878
rect 6006 10850 6034 11103
rect 6342 10962 6370 11159
rect 6342 10929 6370 10934
rect 6006 10817 6034 10822
rect 5334 10767 5335 10793
rect 5361 10767 5362 10793
rect 5334 10761 5362 10767
rect 6398 10794 6426 11438
rect 6510 11130 6538 11495
rect 6510 11097 6538 11102
rect 7014 11746 7042 11751
rect 6790 11073 6818 11079
rect 6790 11047 6791 11073
rect 6817 11047 6818 11073
rect 6790 10962 6818 11047
rect 7014 11018 7042 11718
rect 6818 10934 6874 10962
rect 6790 10929 6818 10934
rect 6398 10761 6426 10766
rect 5670 10738 5698 10743
rect 5670 10691 5698 10710
rect 6734 10737 6762 10743
rect 6734 10711 6735 10737
rect 6761 10711 6762 10737
rect 6734 10682 6762 10711
rect 6734 10649 6762 10654
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 6846 10458 6874 10934
rect 6958 10794 6986 10799
rect 6958 10747 6986 10766
rect 7014 10793 7042 10990
rect 7406 10962 7434 12278
rect 7462 11746 7490 13006
rect 7742 12810 7770 13062
rect 7574 12782 7770 12810
rect 7518 12642 7546 12647
rect 7574 12642 7602 12782
rect 7630 12698 7658 12703
rect 7742 12698 7770 12703
rect 7630 12697 7770 12698
rect 7630 12671 7631 12697
rect 7657 12671 7743 12697
rect 7769 12671 7770 12697
rect 7630 12670 7770 12671
rect 7630 12665 7658 12670
rect 7742 12665 7770 12670
rect 7854 12698 7882 12703
rect 7854 12651 7882 12670
rect 7910 12697 7938 13119
rect 8078 13090 8106 13426
rect 8134 13258 8162 13455
rect 8134 13225 8162 13230
rect 8134 13090 8162 13095
rect 8358 13090 8386 13846
rect 8470 13841 8498 13846
rect 8694 13594 8722 13846
rect 8694 13561 8722 13566
rect 8078 13089 8386 13090
rect 8078 13063 8135 13089
rect 8161 13063 8386 13089
rect 8078 13062 8386 13063
rect 8750 13145 8778 14238
rect 9030 13762 9058 18999
rect 9758 18746 9786 20600
rect 11102 19081 11130 20600
rect 12110 19138 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12110 19105 12138 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 11102 19055 11103 19081
rect 11129 19055 11130 19081
rect 11102 19049 11130 19055
rect 11774 19025 11802 19031
rect 11774 18999 11775 19025
rect 11801 18999 11802 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9758 18713 9786 18718
rect 10374 18746 10402 18751
rect 10374 18699 10402 18718
rect 9870 18634 9898 18639
rect 9478 18633 9898 18634
rect 9478 18607 9871 18633
rect 9897 18607 9898 18633
rect 9478 18606 9898 18607
rect 9366 14266 9394 14271
rect 9366 14219 9394 14238
rect 9478 14266 9506 18606
rect 9870 18601 9898 18606
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9478 14219 9506 14238
rect 9534 14377 9562 14383
rect 9534 14351 9535 14377
rect 9561 14351 9562 14377
rect 9086 13874 9114 13879
rect 9086 13873 9394 13874
rect 9086 13847 9087 13873
rect 9113 13847 9394 13873
rect 9086 13846 9394 13847
rect 9086 13841 9114 13846
rect 9030 13734 9226 13762
rect 9198 13593 9226 13734
rect 9366 13649 9394 13846
rect 9366 13623 9367 13649
rect 9393 13623 9394 13649
rect 9366 13617 9394 13623
rect 9422 13650 9450 13655
rect 9198 13567 9199 13593
rect 9225 13567 9226 13593
rect 8862 13258 8890 13263
rect 8862 13211 8890 13230
rect 9198 13257 9226 13567
rect 9422 13482 9450 13622
rect 9534 13649 9562 14351
rect 10150 14266 10178 14271
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9534 13623 9535 13649
rect 9561 13623 9562 13649
rect 9534 13617 9562 13623
rect 9814 13930 9842 13935
rect 9758 13594 9786 13599
rect 9758 13547 9786 13566
rect 9422 13481 9562 13482
rect 9422 13455 9423 13481
rect 9449 13455 9562 13481
rect 9422 13454 9562 13455
rect 9422 13449 9450 13454
rect 9198 13231 9199 13257
rect 9225 13231 9226 13257
rect 9198 13225 9226 13231
rect 9534 13257 9562 13454
rect 9534 13231 9535 13257
rect 9561 13231 9562 13257
rect 9534 13225 9562 13231
rect 9086 13201 9114 13207
rect 9086 13175 9087 13201
rect 9113 13175 9114 13201
rect 8750 13119 8751 13145
rect 8777 13119 8778 13145
rect 7910 12671 7911 12697
rect 7937 12671 7938 12697
rect 7518 12641 7602 12642
rect 7518 12615 7519 12641
rect 7545 12615 7602 12641
rect 7518 12614 7602 12615
rect 7518 12609 7546 12614
rect 7574 12586 7602 12614
rect 7910 12642 7938 12671
rect 7574 12558 7658 12586
rect 7462 11713 7490 11718
rect 7574 11634 7602 11639
rect 7574 11587 7602 11606
rect 7406 10929 7434 10934
rect 7518 11522 7546 11527
rect 7350 10906 7378 10911
rect 7350 10859 7378 10878
rect 7182 10850 7210 10855
rect 7182 10803 7210 10822
rect 7014 10767 7015 10793
rect 7041 10767 7042 10793
rect 7014 10761 7042 10767
rect 7294 10794 7322 10799
rect 6790 10430 6846 10458
rect 4998 10010 5026 10015
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 966 9673 994 9679
rect 966 9647 967 9673
rect 993 9647 994 9673
rect 966 9450 994 9647
rect 4998 9674 5026 9982
rect 4998 9627 5026 9646
rect 2142 9618 2170 9623
rect 2142 9571 2170 9590
rect 6454 9618 6482 9623
rect 6454 9571 6482 9590
rect 6790 9618 6818 10430
rect 6846 10411 6874 10430
rect 7182 10402 7210 10407
rect 7294 10402 7322 10766
rect 7182 10401 7322 10402
rect 7182 10375 7183 10401
rect 7209 10375 7322 10401
rect 7182 10374 7322 10375
rect 7406 10793 7434 10799
rect 7406 10767 7407 10793
rect 7433 10767 7434 10793
rect 7182 10369 7210 10374
rect 7014 10345 7042 10351
rect 7014 10319 7015 10345
rect 7041 10319 7042 10345
rect 7014 10094 7042 10319
rect 7070 10289 7098 10295
rect 7070 10263 7071 10289
rect 7097 10263 7098 10289
rect 7070 10178 7098 10263
rect 7294 10289 7322 10295
rect 7294 10263 7295 10289
rect 7321 10263 7322 10289
rect 7294 10178 7322 10263
rect 7070 10150 7322 10178
rect 7014 10066 7210 10094
rect 7126 10010 7154 10015
rect 7126 9963 7154 9982
rect 966 9417 994 9422
rect 6062 9561 6090 9567
rect 6062 9535 6063 9561
rect 6089 9535 6090 9561
rect 6062 9338 6090 9535
rect 6062 9305 6090 9310
rect 6734 9562 6762 9567
rect 6734 9225 6762 9534
rect 6734 9199 6735 9225
rect 6761 9199 6762 9225
rect 6734 9193 6762 9199
rect 6790 9505 6818 9590
rect 7182 9617 7210 10066
rect 7182 9591 7183 9617
rect 7209 9591 7210 9617
rect 6790 9479 6791 9505
rect 6817 9479 6818 9505
rect 6678 9169 6706 9175
rect 6678 9143 6679 9169
rect 6705 9143 6706 9169
rect 6678 9114 6706 9143
rect 6678 9081 6706 9086
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 5838 8498 5866 8503
rect 5838 8451 5866 8470
rect 5502 8442 5530 8447
rect 5502 8395 5530 8414
rect 6342 8386 6370 8391
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 6342 7657 6370 8358
rect 6790 8386 6818 9479
rect 7126 9562 7154 9567
rect 7126 9450 7154 9534
rect 7070 9422 7154 9450
rect 6958 9226 6986 9231
rect 6958 9179 6986 9198
rect 6902 9170 6930 9175
rect 6902 9123 6930 9142
rect 7070 8833 7098 9422
rect 7126 9338 7154 9343
rect 7126 9291 7154 9310
rect 7182 9058 7210 9591
rect 7238 9898 7266 9903
rect 7294 9898 7322 10150
rect 7406 10234 7434 10767
rect 7238 9897 7322 9898
rect 7238 9871 7239 9897
rect 7265 9871 7322 9897
rect 7238 9870 7322 9871
rect 7350 10121 7378 10127
rect 7350 10095 7351 10121
rect 7377 10095 7378 10121
rect 7238 9618 7266 9870
rect 7350 9730 7378 10095
rect 7406 10094 7434 10206
rect 7462 10289 7490 10295
rect 7462 10263 7463 10289
rect 7489 10263 7490 10289
rect 7462 10178 7490 10263
rect 7462 10145 7490 10150
rect 7406 10066 7490 10094
rect 7406 10009 7434 10015
rect 7406 9983 7407 10009
rect 7433 9983 7434 10009
rect 7406 9898 7434 9983
rect 7462 9954 7490 10066
rect 7518 10065 7546 11494
rect 7574 10794 7602 10799
rect 7574 10747 7602 10766
rect 7518 10039 7519 10065
rect 7545 10039 7546 10065
rect 7518 10033 7546 10039
rect 7462 9926 7574 9954
rect 7406 9865 7434 9870
rect 7546 9786 7574 9926
rect 7238 9585 7266 9590
rect 7294 9702 7378 9730
rect 7406 9758 7574 9786
rect 7238 9505 7266 9511
rect 7238 9479 7239 9505
rect 7265 9479 7266 9505
rect 7238 9225 7266 9479
rect 7238 9199 7239 9225
rect 7265 9199 7266 9225
rect 7238 9193 7266 9199
rect 7294 9225 7322 9702
rect 7294 9199 7295 9225
rect 7321 9199 7322 9225
rect 7294 9193 7322 9199
rect 7350 9561 7378 9567
rect 7350 9535 7351 9561
rect 7377 9535 7378 9561
rect 7350 9506 7378 9535
rect 7182 9025 7210 9030
rect 7238 9114 7266 9119
rect 7070 8807 7071 8833
rect 7097 8807 7098 8833
rect 7070 8801 7098 8807
rect 6958 8721 6986 8727
rect 6958 8695 6959 8721
rect 6985 8695 6986 8721
rect 6958 8498 6986 8695
rect 7238 8553 7266 9086
rect 7350 8889 7378 9478
rect 7406 9281 7434 9758
rect 7630 9730 7658 12558
rect 7910 11970 7938 12614
rect 7910 11937 7938 11942
rect 8134 12362 8162 13062
rect 8078 11858 8106 11863
rect 8134 11858 8162 12334
rect 8106 11830 8162 11858
rect 8190 12810 8218 12815
rect 8190 12641 8218 12782
rect 8190 12615 8191 12641
rect 8217 12615 8218 12641
rect 7910 11578 7938 11583
rect 8078 11578 8106 11830
rect 8190 11746 8218 12615
rect 8750 12306 8778 13119
rect 8806 13145 8834 13151
rect 8806 13119 8807 13145
rect 8833 13119 8834 13145
rect 8806 13090 8834 13119
rect 9030 13146 9058 13151
rect 9086 13146 9114 13175
rect 9030 13145 9114 13146
rect 9030 13119 9031 13145
rect 9057 13119 9114 13145
rect 9030 13118 9114 13119
rect 9254 13145 9282 13151
rect 9254 13119 9255 13145
rect 9281 13119 9282 13145
rect 9030 13113 9058 13118
rect 8806 13057 8834 13062
rect 9254 12642 9282 13119
rect 9646 13146 9674 13151
rect 9814 13146 9842 13902
rect 10150 13873 10178 14238
rect 10150 13847 10151 13873
rect 10177 13847 10178 13873
rect 10150 13841 10178 13847
rect 10654 13930 10682 13935
rect 10262 13706 10290 13711
rect 10150 13481 10178 13487
rect 10150 13455 10151 13481
rect 10177 13455 10178 13481
rect 10150 13426 10178 13455
rect 10150 13393 10178 13398
rect 10206 13481 10234 13487
rect 10206 13455 10207 13481
rect 10233 13455 10234 13481
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9870 13146 9898 13151
rect 9814 13145 9898 13146
rect 9814 13119 9871 13145
rect 9897 13119 9898 13145
rect 9814 13118 9898 13119
rect 9646 13099 9674 13118
rect 9870 13113 9898 13118
rect 9254 12609 9282 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10206 12474 10234 13455
rect 10262 13481 10290 13678
rect 10374 13650 10402 13655
rect 10374 13537 10402 13622
rect 10374 13511 10375 13537
rect 10401 13511 10402 13537
rect 10374 13505 10402 13511
rect 10262 13455 10263 13481
rect 10289 13455 10290 13481
rect 10262 13449 10290 13455
rect 10654 13482 10682 13902
rect 11046 13873 11074 13879
rect 11046 13847 11047 13873
rect 11073 13847 11074 13873
rect 11046 13594 11074 13847
rect 11718 13874 11746 13879
rect 11438 13706 11466 13711
rect 11270 13650 11298 13655
rect 11102 13594 11130 13599
rect 11046 13593 11130 13594
rect 11046 13567 11103 13593
rect 11129 13567 11130 13593
rect 11046 13566 11130 13567
rect 11102 13561 11130 13566
rect 11158 13594 11186 13599
rect 10934 13537 10962 13543
rect 10934 13511 10935 13537
rect 10961 13511 10962 13537
rect 10654 13449 10682 13454
rect 10878 13482 10906 13487
rect 10934 13482 10962 13511
rect 10934 13454 11018 13482
rect 10318 13425 10346 13431
rect 10318 13399 10319 13425
rect 10345 13399 10346 13425
rect 10262 13202 10290 13207
rect 10318 13202 10346 13399
rect 10878 13370 10906 13454
rect 10878 13342 10962 13370
rect 10262 13201 10346 13202
rect 10262 13175 10263 13201
rect 10289 13175 10346 13201
rect 10262 13174 10346 13175
rect 10262 13169 10290 13174
rect 10206 12446 10458 12474
rect 9590 12418 9618 12423
rect 9590 12371 9618 12390
rect 9758 12361 9786 12367
rect 9758 12335 9759 12361
rect 9785 12335 9786 12361
rect 8750 12278 8946 12306
rect 8470 11969 8498 11975
rect 8470 11943 8471 11969
rect 8497 11943 8498 11969
rect 8470 11858 8498 11943
rect 8470 11825 8498 11830
rect 8862 11913 8890 11919
rect 8862 11887 8863 11913
rect 8889 11887 8890 11913
rect 8190 11713 8218 11718
rect 8694 11746 8722 11751
rect 8190 11634 8218 11639
rect 8190 11587 8218 11606
rect 7910 11577 8106 11578
rect 7910 11551 7911 11577
rect 7937 11551 8106 11577
rect 7910 11550 8106 11551
rect 8134 11577 8162 11583
rect 8134 11551 8135 11577
rect 8161 11551 8162 11577
rect 7798 11186 7826 11191
rect 7798 10849 7826 11158
rect 7910 10962 7938 11550
rect 7910 10929 7938 10934
rect 8078 11186 8106 11191
rect 8078 10962 8106 11158
rect 8078 10929 8106 10934
rect 7798 10823 7799 10849
rect 7825 10823 7826 10849
rect 7686 10738 7714 10743
rect 7686 10691 7714 10710
rect 7742 10458 7770 10463
rect 7742 10411 7770 10430
rect 7574 9702 7658 9730
rect 7406 9255 7407 9281
rect 7433 9255 7434 9281
rect 7406 9249 7434 9255
rect 7462 9674 7490 9679
rect 7462 9561 7490 9646
rect 7574 9673 7602 9702
rect 7574 9647 7575 9673
rect 7601 9647 7602 9673
rect 7574 9641 7602 9647
rect 7630 9618 7658 9623
rect 7630 9571 7658 9590
rect 7462 9535 7463 9561
rect 7489 9535 7490 9561
rect 7350 8863 7351 8889
rect 7377 8863 7378 8889
rect 7350 8857 7378 8863
rect 7462 9226 7490 9535
rect 7742 9562 7770 9567
rect 7742 9515 7770 9534
rect 7518 9282 7546 9287
rect 7518 9235 7546 9254
rect 7462 8834 7490 9198
rect 7742 8834 7770 8839
rect 7462 8833 7770 8834
rect 7462 8807 7743 8833
rect 7769 8807 7770 8833
rect 7462 8806 7770 8807
rect 7742 8801 7770 8806
rect 7238 8527 7239 8553
rect 7265 8527 7266 8553
rect 7238 8521 7266 8527
rect 7574 8721 7602 8727
rect 7798 8722 7826 10823
rect 8078 10849 8106 10855
rect 8078 10823 8079 10849
rect 8105 10823 8106 10849
rect 7910 10793 7938 10799
rect 7910 10767 7911 10793
rect 7937 10767 7938 10793
rect 7910 10738 7938 10767
rect 7910 10705 7938 10710
rect 8022 10794 8050 10799
rect 8022 10122 8050 10766
rect 8078 10234 8106 10823
rect 8134 10737 8162 11551
rect 8246 11577 8274 11583
rect 8246 11551 8247 11577
rect 8273 11551 8274 11577
rect 8190 11298 8218 11303
rect 8246 11298 8274 11551
rect 8414 11578 8442 11583
rect 8414 11531 8442 11550
rect 8190 11297 8274 11298
rect 8190 11271 8191 11297
rect 8217 11271 8274 11297
rect 8190 11270 8274 11271
rect 8190 11265 8218 11270
rect 8694 11242 8722 11718
rect 8806 11690 8834 11695
rect 8862 11690 8890 11887
rect 8806 11689 8890 11690
rect 8806 11663 8807 11689
rect 8833 11663 8890 11689
rect 8806 11662 8890 11663
rect 8806 11657 8834 11662
rect 8190 11130 8218 11135
rect 8190 11083 8218 11102
rect 8246 11130 8274 11135
rect 8246 11129 8386 11130
rect 8246 11103 8247 11129
rect 8273 11103 8386 11129
rect 8246 11102 8386 11103
rect 8246 11097 8274 11102
rect 8246 10962 8274 10967
rect 8134 10711 8135 10737
rect 8161 10711 8162 10737
rect 8134 10705 8162 10711
rect 8190 10793 8218 10799
rect 8190 10767 8191 10793
rect 8217 10767 8218 10793
rect 8078 10201 8106 10206
rect 8078 10122 8106 10127
rect 8190 10122 8218 10767
rect 8022 10121 8106 10122
rect 8022 10095 8079 10121
rect 8105 10095 8106 10121
rect 8022 10094 8106 10095
rect 8078 10089 8106 10094
rect 8134 10094 8190 10122
rect 7966 10066 7994 10071
rect 7966 10009 7994 10038
rect 7966 9983 7967 10009
rect 7993 9983 7994 10009
rect 7966 9618 7994 9983
rect 8134 9674 8162 10094
rect 8190 10089 8218 10094
rect 8246 10121 8274 10934
rect 8302 10794 8330 10799
rect 8302 10747 8330 10766
rect 8246 10095 8247 10121
rect 8273 10095 8274 10121
rect 8246 10089 8274 10095
rect 8358 10094 8386 11102
rect 8470 11129 8498 11135
rect 8470 11103 8471 11129
rect 8497 11103 8498 11129
rect 7966 9585 7994 9590
rect 8022 9646 8162 9674
rect 8302 10066 8386 10094
rect 8414 11073 8442 11079
rect 8414 11047 8415 11073
rect 8441 11047 8442 11073
rect 8414 10066 8442 11047
rect 8470 10682 8498 11103
rect 8694 10794 8722 11214
rect 8750 11577 8778 11583
rect 8750 11551 8751 11577
rect 8777 11551 8778 11577
rect 8750 11186 8778 11551
rect 8862 11578 8890 11583
rect 8918 11578 8946 12278
rect 9758 12250 9786 12335
rect 10206 12362 10234 12367
rect 10206 12315 10234 12334
rect 9982 12305 10010 12311
rect 9982 12279 9983 12305
rect 10009 12279 10010 12305
rect 9926 12250 9954 12255
rect 9758 12249 9954 12250
rect 9758 12223 9927 12249
rect 9953 12223 9954 12249
rect 9758 12222 9954 12223
rect 8890 11550 8946 11578
rect 8974 11633 9002 11639
rect 8974 11607 8975 11633
rect 9001 11607 9002 11633
rect 8862 11531 8890 11550
rect 8750 11153 8778 11158
rect 8694 10761 8722 10766
rect 8862 10793 8890 10799
rect 8862 10767 8863 10793
rect 8889 10767 8890 10793
rect 8470 10649 8498 10654
rect 8862 10682 8890 10767
rect 8862 10649 8890 10654
rect 8974 10346 9002 11607
rect 9254 11633 9282 11639
rect 9254 11607 9255 11633
rect 9281 11607 9282 11633
rect 9254 11578 9282 11607
rect 9422 11634 9450 11639
rect 9758 11634 9786 12222
rect 9926 12217 9954 12222
rect 9926 12026 9954 12031
rect 9982 12026 10010 12279
rect 9926 12025 10234 12026
rect 9926 11999 9927 12025
rect 9953 11999 10234 12025
rect 9926 11998 10234 11999
rect 9926 11993 9954 11998
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10150 11689 10178 11998
rect 10206 11969 10234 11998
rect 10206 11943 10207 11969
rect 10233 11943 10234 11969
rect 10206 11937 10234 11943
rect 10150 11663 10151 11689
rect 10177 11663 10178 11689
rect 10150 11657 10178 11663
rect 10374 11857 10402 11863
rect 10374 11831 10375 11857
rect 10401 11831 10402 11857
rect 10374 11746 10402 11831
rect 10038 11634 10066 11639
rect 9422 11633 9842 11634
rect 9422 11607 9423 11633
rect 9449 11607 9842 11633
rect 9422 11606 9842 11607
rect 9422 11601 9450 11606
rect 9254 11545 9282 11550
rect 9814 11577 9842 11606
rect 9814 11551 9815 11577
rect 9841 11551 9842 11577
rect 9814 11545 9842 11551
rect 9590 11522 9618 11527
rect 9590 11475 9618 11494
rect 9310 11186 9338 11191
rect 9030 11130 9058 11135
rect 9030 10905 9058 11102
rect 9086 11074 9114 11079
rect 9086 11027 9114 11046
rect 9254 11074 9282 11079
rect 9310 11074 9338 11158
rect 9646 11185 9674 11191
rect 9646 11159 9647 11185
rect 9673 11159 9674 11185
rect 9422 11130 9450 11135
rect 9422 11083 9450 11102
rect 9590 11129 9618 11135
rect 9590 11103 9591 11129
rect 9617 11103 9618 11129
rect 9254 11073 9338 11074
rect 9254 11047 9255 11073
rect 9281 11047 9338 11073
rect 9254 11046 9338 11047
rect 9254 11041 9282 11046
rect 9030 10879 9031 10905
rect 9057 10879 9058 10905
rect 9030 10873 9058 10879
rect 9198 10794 9226 10799
rect 8862 10318 9002 10346
rect 9030 10766 9198 10794
rect 7574 8695 7575 8721
rect 7601 8695 7602 8721
rect 6958 8465 6986 8470
rect 7574 8498 7602 8695
rect 7686 8694 7826 8722
rect 7854 9169 7882 9175
rect 7854 9143 7855 9169
rect 7881 9143 7882 9169
rect 7854 8722 7882 9143
rect 8022 9058 8050 9646
rect 8134 9562 8162 9567
rect 8302 9562 8330 10066
rect 8414 10033 8442 10038
rect 8526 10234 8554 10239
rect 8134 9561 8218 9562
rect 8134 9535 8135 9561
rect 8161 9535 8218 9561
rect 8134 9534 8218 9535
rect 8134 9529 8162 9534
rect 8134 9226 8162 9231
rect 8078 9114 8106 9119
rect 8134 9114 8162 9198
rect 8106 9086 8162 9114
rect 8078 9081 8106 9086
rect 7910 9030 8050 9058
rect 7910 8777 7938 9030
rect 7910 8751 7911 8777
rect 7937 8751 7938 8777
rect 7910 8745 7938 8751
rect 7966 8946 7994 8951
rect 7630 8498 7658 8503
rect 7574 8497 7658 8498
rect 7574 8471 7631 8497
rect 7657 8471 7658 8497
rect 7574 8470 7658 8471
rect 6790 8353 6818 8358
rect 6902 8442 6930 8447
rect 6902 8385 6930 8414
rect 7350 8442 7378 8447
rect 7350 8395 7378 8414
rect 7574 8442 7602 8470
rect 7630 8465 7658 8470
rect 7574 8409 7602 8414
rect 6902 8359 6903 8385
rect 6929 8359 6930 8385
rect 6902 8353 6930 8359
rect 7630 8386 7658 8391
rect 7630 7993 7658 8358
rect 7686 8162 7714 8694
rect 7854 8498 7882 8694
rect 7910 8554 7938 8559
rect 7966 8554 7994 8918
rect 8134 8889 8162 9086
rect 8190 9169 8218 9534
rect 8302 9529 8330 9534
rect 8358 10010 8386 10015
rect 8190 9143 8191 9169
rect 8217 9143 8218 9169
rect 8190 9114 8218 9143
rect 8190 9081 8218 9086
rect 8246 9170 8274 9175
rect 8134 8863 8135 8889
rect 8161 8863 8162 8889
rect 8134 8857 8162 8863
rect 8246 8945 8274 9142
rect 8358 9114 8386 9982
rect 8414 9617 8442 9623
rect 8414 9591 8415 9617
rect 8441 9591 8442 9617
rect 8414 9226 8442 9591
rect 8526 9618 8554 10206
rect 8862 9730 8890 10318
rect 8974 9954 9002 9959
rect 8862 9683 8890 9702
rect 8918 9926 8974 9954
rect 8526 9590 8722 9618
rect 8526 9561 8554 9590
rect 8526 9535 8527 9561
rect 8553 9535 8554 9561
rect 8526 9529 8554 9535
rect 8694 9561 8722 9590
rect 8694 9535 8695 9561
rect 8721 9535 8722 9561
rect 8694 9529 8722 9535
rect 8918 9561 8946 9926
rect 8974 9907 9002 9926
rect 8918 9535 8919 9561
rect 8945 9535 8946 9561
rect 8806 9505 8834 9511
rect 8806 9479 8807 9505
rect 8833 9479 8834 9505
rect 8414 9193 8442 9198
rect 8694 9225 8722 9231
rect 8694 9199 8695 9225
rect 8721 9199 8722 9225
rect 8358 9086 8442 9114
rect 8246 8919 8247 8945
rect 8273 8919 8274 8945
rect 7910 8553 7994 8554
rect 7910 8527 7911 8553
rect 7937 8527 7994 8553
rect 7910 8526 7994 8527
rect 8246 8834 8274 8919
rect 8414 8945 8442 9086
rect 8414 8919 8415 8945
rect 8441 8919 8442 8945
rect 8414 8913 8442 8919
rect 8246 8553 8274 8806
rect 8582 8834 8610 8839
rect 8694 8834 8722 9199
rect 8610 8806 8722 8834
rect 8582 8787 8610 8806
rect 8750 8778 8778 8783
rect 8806 8778 8834 9479
rect 8918 9282 8946 9535
rect 8918 9249 8946 9254
rect 8974 9226 9002 9231
rect 8974 9179 9002 9198
rect 8750 8777 8834 8778
rect 8750 8751 8751 8777
rect 8777 8751 8834 8777
rect 8750 8750 8834 8751
rect 8750 8745 8778 8750
rect 8246 8527 8247 8553
rect 8273 8527 8274 8553
rect 7910 8521 7938 8526
rect 8246 8521 8274 8527
rect 8806 8554 8834 8750
rect 8806 8521 8834 8526
rect 7798 8470 7882 8498
rect 7798 8442 7826 8470
rect 8078 8442 8106 8447
rect 7798 8409 7826 8414
rect 7854 8441 8106 8442
rect 7854 8415 8079 8441
rect 8105 8415 8106 8441
rect 7854 8414 8106 8415
rect 7742 8330 7770 8335
rect 7854 8330 7882 8414
rect 8078 8409 8106 8414
rect 9030 8442 9058 10766
rect 9198 10747 9226 10766
rect 9254 10738 9282 10743
rect 9254 10691 9282 10710
rect 9142 10346 9170 10351
rect 9310 10346 9338 11046
rect 9534 11074 9562 11079
rect 9534 10793 9562 11046
rect 9590 11018 9618 11103
rect 9590 10985 9618 10990
rect 9534 10767 9535 10793
rect 9561 10767 9562 10793
rect 9534 10761 9562 10767
rect 9142 9953 9170 10318
rect 9142 9927 9143 9953
rect 9169 9927 9170 9953
rect 9142 9921 9170 9927
rect 9198 10318 9338 10346
rect 9366 10682 9394 10687
rect 9646 10682 9674 11159
rect 9926 11185 9954 11191
rect 9926 11159 9927 11185
rect 9953 11159 9954 11185
rect 9926 11074 9954 11159
rect 10038 11074 10066 11606
rect 10318 11634 10346 11639
rect 10318 11587 10346 11606
rect 10094 11578 10122 11583
rect 10094 11186 10122 11550
rect 10094 11139 10122 11158
rect 9926 11046 10122 11074
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9366 10681 9674 10682
rect 9366 10655 9367 10681
rect 9393 10655 9674 10681
rect 9366 10654 9674 10655
rect 9198 10009 9226 10318
rect 9198 9983 9199 10009
rect 9225 9983 9226 10009
rect 9086 9618 9114 9623
rect 9086 9571 9114 9590
rect 9198 9618 9226 9983
rect 9198 9585 9226 9590
rect 9254 10234 9282 10239
rect 9254 9562 9282 10206
rect 9366 10010 9394 10654
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10038 10122 10066 10127
rect 10038 10075 10066 10094
rect 9590 10066 9618 10071
rect 9814 10066 9842 10071
rect 9366 9977 9394 9982
rect 9534 10009 9562 10015
rect 9534 9983 9535 10009
rect 9561 9983 9562 10009
rect 9534 9954 9562 9983
rect 9534 9921 9562 9926
rect 9422 9562 9450 9567
rect 9254 9561 9394 9562
rect 9254 9535 9255 9561
rect 9281 9535 9394 9561
rect 9254 9534 9394 9535
rect 9254 9529 9282 9534
rect 9310 8554 9338 8559
rect 9310 8507 9338 8526
rect 9254 8498 9282 8503
rect 9254 8442 9282 8470
rect 9254 8414 9338 8442
rect 7742 8329 7882 8330
rect 7742 8303 7743 8329
rect 7769 8303 7882 8329
rect 7742 8302 7882 8303
rect 7742 8297 7770 8302
rect 7742 8162 7770 8167
rect 7686 8134 7742 8162
rect 7742 8115 7770 8134
rect 7630 7967 7631 7993
rect 7657 7967 7658 7993
rect 7630 7961 7658 7967
rect 6678 7938 6706 7943
rect 6678 7713 6706 7910
rect 6678 7687 6679 7713
rect 6705 7687 6706 7713
rect 6678 7681 6706 7687
rect 7014 7937 7042 7943
rect 7014 7911 7015 7937
rect 7041 7911 7042 7937
rect 6342 7631 6343 7657
rect 6369 7631 6370 7657
rect 6342 7602 6370 7631
rect 6342 7569 6370 7574
rect 7014 7602 7042 7911
rect 7686 7938 7714 7943
rect 7686 7891 7714 7910
rect 7686 7714 7714 7719
rect 7014 7569 7042 7574
rect 7350 7602 7378 7607
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7350 7265 7378 7574
rect 7686 7321 7714 7686
rect 7742 7602 7770 7607
rect 7798 7602 7826 8302
rect 8694 8162 8722 8167
rect 8694 8049 8722 8134
rect 8694 8023 8695 8049
rect 8721 8023 8722 8049
rect 8694 8017 8722 8023
rect 9030 8049 9058 8414
rect 9254 8329 9282 8335
rect 9254 8303 9255 8329
rect 9281 8303 9282 8329
rect 9030 8023 9031 8049
rect 9057 8023 9058 8049
rect 9030 8017 9058 8023
rect 9086 8105 9114 8111
rect 9086 8079 9087 8105
rect 9113 8079 9114 8105
rect 8806 7994 8834 7999
rect 8806 7947 8834 7966
rect 8862 7993 8890 7999
rect 8862 7967 8863 7993
rect 8889 7967 8890 7993
rect 7742 7601 7826 7602
rect 7742 7575 7743 7601
rect 7769 7575 7826 7601
rect 7742 7574 7826 7575
rect 7966 7602 7994 7621
rect 7742 7569 7770 7574
rect 7966 7569 7994 7574
rect 8750 7602 8778 7621
rect 8750 7546 8834 7574
rect 7686 7295 7687 7321
rect 7713 7295 7714 7321
rect 7686 7289 7714 7295
rect 8750 7322 8778 7327
rect 8750 7275 8778 7294
rect 7350 7239 7351 7265
rect 7377 7239 7378 7265
rect 7350 7233 7378 7239
rect 8806 7266 8834 7546
rect 8862 7378 8890 7967
rect 9086 7713 9114 8079
rect 9086 7687 9087 7713
rect 9113 7687 9114 7713
rect 9086 7681 9114 7687
rect 9142 7714 9170 7719
rect 9142 7667 9170 7686
rect 9254 7713 9282 8303
rect 9310 8161 9338 8414
rect 9310 8135 9311 8161
rect 9337 8135 9338 8161
rect 9310 8129 9338 8135
rect 9366 8162 9394 9534
rect 9422 8553 9450 9534
rect 9590 8554 9618 10038
rect 9758 10038 9814 10066
rect 9758 9506 9786 10038
rect 9814 10019 9842 10038
rect 9982 10010 10010 10015
rect 9982 9618 10010 9982
rect 9758 9473 9786 9478
rect 9814 9617 10010 9618
rect 9814 9591 9983 9617
rect 10009 9591 10010 9617
rect 9814 9590 10010 9591
rect 9814 9226 9842 9590
rect 9982 9585 10010 9590
rect 10038 9506 10066 9525
rect 10038 9473 10066 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9814 9193 9842 9198
rect 10094 9225 10122 11046
rect 10374 10962 10402 11718
rect 10430 11242 10458 12446
rect 10934 12361 10962 13342
rect 10934 12335 10935 12361
rect 10961 12335 10962 12361
rect 10934 12329 10962 12335
rect 10990 12082 11018 13454
rect 11102 13481 11130 13487
rect 11102 13455 11103 13481
rect 11129 13455 11130 13481
rect 11102 13426 11130 13455
rect 11158 13481 11186 13566
rect 11158 13455 11159 13481
rect 11185 13455 11186 13481
rect 11158 13449 11186 13455
rect 11270 13537 11298 13622
rect 11270 13511 11271 13537
rect 11297 13511 11298 13537
rect 11102 12194 11130 13398
rect 11270 12866 11298 13511
rect 11438 13481 11466 13678
rect 11662 13594 11690 13599
rect 11662 13547 11690 13566
rect 11718 13593 11746 13846
rect 11718 13567 11719 13593
rect 11745 13567 11746 13593
rect 11718 13561 11746 13567
rect 11438 13455 11439 13481
rect 11465 13455 11466 13481
rect 11438 13449 11466 13455
rect 11494 13510 11634 13538
rect 11494 13481 11522 13510
rect 11494 13455 11495 13481
rect 11521 13455 11522 13481
rect 11326 13090 11354 13095
rect 11494 13090 11522 13455
rect 11606 13482 11634 13510
rect 11774 13482 11802 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 12110 15946 12306 15974
rect 12110 13874 12138 15946
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 12110 13827 12138 13846
rect 12390 13873 12418 13879
rect 12390 13847 12391 13873
rect 12417 13847 12418 13873
rect 11606 13454 11802 13482
rect 12054 13482 12082 13487
rect 11550 13426 11578 13431
rect 11550 13257 11578 13398
rect 11550 13231 11551 13257
rect 11577 13231 11578 13257
rect 11550 13225 11578 13231
rect 11326 13089 11522 13090
rect 11326 13063 11327 13089
rect 11353 13063 11522 13089
rect 11326 13062 11522 13063
rect 11326 13057 11354 13062
rect 11326 12866 11354 12871
rect 11270 12865 11354 12866
rect 11270 12839 11327 12865
rect 11353 12839 11354 12865
rect 11270 12838 11354 12839
rect 11326 12833 11354 12838
rect 11494 12810 11522 12815
rect 11494 12753 11522 12782
rect 11494 12727 11495 12753
rect 11521 12727 11522 12753
rect 11494 12721 11522 12727
rect 12054 12753 12082 13454
rect 12390 13482 12418 13847
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 12418 13454 12474 13482
rect 12390 13449 12418 13454
rect 12054 12727 12055 12753
rect 12081 12727 12082 12753
rect 12054 12721 12082 12727
rect 11606 12698 11634 12703
rect 11606 12651 11634 12670
rect 12390 12698 12418 12703
rect 12390 12651 12418 12670
rect 11550 12642 11578 12647
rect 11270 12306 11298 12311
rect 11270 12305 11410 12306
rect 11270 12279 11271 12305
rect 11297 12279 11410 12305
rect 11270 12278 11410 12279
rect 11270 12273 11298 12278
rect 11102 12166 11242 12194
rect 10990 12054 11130 12082
rect 10654 11970 10682 11975
rect 10654 11913 10682 11942
rect 10654 11887 10655 11913
rect 10681 11887 10682 11913
rect 10654 11881 10682 11887
rect 10766 11969 10794 11975
rect 11046 11970 11074 11975
rect 10766 11943 10767 11969
rect 10793 11943 10794 11969
rect 10766 11746 10794 11943
rect 10878 11969 11074 11970
rect 10878 11943 11047 11969
rect 11073 11943 11074 11969
rect 10878 11942 11074 11943
rect 10766 11713 10794 11718
rect 10822 11802 10850 11807
rect 10822 11633 10850 11774
rect 10822 11607 10823 11633
rect 10849 11607 10850 11633
rect 10654 11578 10682 11583
rect 10654 11531 10682 11550
rect 10766 11410 10794 11415
rect 10598 11242 10626 11247
rect 10430 11241 10626 11242
rect 10430 11215 10599 11241
rect 10625 11215 10626 11241
rect 10430 11214 10626 11215
rect 10598 11209 10626 11214
rect 10766 11185 10794 11382
rect 10766 11159 10767 11185
rect 10793 11159 10794 11185
rect 10766 11153 10794 11159
rect 10374 10929 10402 10934
rect 10654 11129 10682 11135
rect 10654 11103 10655 11129
rect 10681 11103 10682 11129
rect 10206 10570 10234 10575
rect 10150 9618 10178 9623
rect 10206 9618 10234 10542
rect 10654 10290 10682 11103
rect 10766 10962 10794 10967
rect 10766 10401 10794 10934
rect 10766 10375 10767 10401
rect 10793 10375 10794 10401
rect 10766 10346 10794 10375
rect 10766 10313 10794 10318
rect 10654 10257 10682 10262
rect 10262 10010 10290 10015
rect 10262 9963 10290 9982
rect 10822 9954 10850 11607
rect 10878 11186 10906 11942
rect 11046 11937 11074 11942
rect 10878 11139 10906 11158
rect 10934 11185 10962 11191
rect 10934 11159 10935 11185
rect 10961 11159 10962 11185
rect 10934 10906 10962 11159
rect 10934 10570 10962 10878
rect 10934 10537 10962 10542
rect 10990 10402 11018 10407
rect 10990 10401 11074 10402
rect 10990 10375 10991 10401
rect 11017 10375 11074 10401
rect 10990 10374 11074 10375
rect 10990 10369 11018 10374
rect 10878 10066 10906 10071
rect 10990 10066 11018 10071
rect 10906 10065 11018 10066
rect 10906 10039 10991 10065
rect 11017 10039 11018 10065
rect 10906 10038 11018 10039
rect 10878 10033 10906 10038
rect 10990 10033 11018 10038
rect 11046 9954 11074 10374
rect 11102 10122 11130 12054
rect 11158 11970 11186 11975
rect 11158 11923 11186 11942
rect 11214 11690 11242 12166
rect 11270 12138 11298 12143
rect 11270 11969 11298 12110
rect 11382 12025 11410 12278
rect 11550 12138 11578 12614
rect 11550 12105 11578 12110
rect 11662 12641 11690 12647
rect 11662 12615 11663 12641
rect 11689 12615 11690 12641
rect 11662 12026 11690 12615
rect 11998 12418 12026 12423
rect 11382 11999 11383 12025
rect 11409 11999 11410 12025
rect 11382 11993 11410 11999
rect 11438 11998 11690 12026
rect 11886 12362 11914 12367
rect 11270 11943 11271 11969
rect 11297 11943 11298 11969
rect 11270 11802 11298 11943
rect 11270 11769 11298 11774
rect 11382 11914 11410 11919
rect 11438 11914 11466 11998
rect 11382 11913 11466 11914
rect 11382 11887 11383 11913
rect 11409 11887 11466 11913
rect 11382 11886 11466 11887
rect 11718 11969 11746 11975
rect 11718 11943 11719 11969
rect 11745 11943 11746 11969
rect 11214 11662 11354 11690
rect 11158 11129 11186 11135
rect 11158 11103 11159 11129
rect 11185 11103 11186 11129
rect 11158 10962 11186 11103
rect 11158 10929 11186 10934
rect 11270 11129 11298 11135
rect 11270 11103 11271 11129
rect 11297 11103 11298 11129
rect 11102 10089 11130 10094
rect 11214 10345 11242 10351
rect 11214 10319 11215 10345
rect 11241 10319 11242 10345
rect 11214 10010 11242 10319
rect 11214 9977 11242 9982
rect 10822 9926 10906 9954
rect 10150 9617 10234 9618
rect 10150 9591 10151 9617
rect 10177 9591 10234 9617
rect 10150 9590 10234 9591
rect 10654 9618 10682 9623
rect 10150 9585 10178 9590
rect 10654 9571 10682 9590
rect 10822 9562 10850 9567
rect 10822 9515 10850 9534
rect 10766 9338 10794 9343
rect 10094 9199 10095 9225
rect 10121 9199 10122 9225
rect 10094 9170 10122 9199
rect 10094 9137 10122 9142
rect 10206 9281 10234 9287
rect 10206 9255 10207 9281
rect 10233 9255 10234 9281
rect 10206 9058 10234 9255
rect 10150 9030 10206 9058
rect 9702 8834 9730 8839
rect 9422 8527 9423 8553
rect 9449 8527 9450 8553
rect 9422 8521 9450 8527
rect 9478 8526 9618 8554
rect 9646 8806 9702 8834
rect 9366 8129 9394 8134
rect 9422 8162 9450 8167
rect 9478 8162 9506 8526
rect 9590 8442 9618 8447
rect 9646 8442 9674 8806
rect 9702 8801 9730 8806
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9926 8554 9954 8559
rect 9814 8498 9842 8503
rect 9814 8451 9842 8470
rect 9926 8497 9954 8526
rect 9926 8471 9927 8497
rect 9953 8471 9954 8497
rect 9590 8441 9674 8442
rect 9590 8415 9591 8441
rect 9617 8415 9674 8441
rect 9590 8414 9674 8415
rect 9590 8409 9618 8414
rect 9590 8330 9618 8335
rect 9422 8161 9506 8162
rect 9422 8135 9423 8161
rect 9449 8135 9506 8161
rect 9422 8134 9506 8135
rect 9422 8129 9450 8134
rect 9254 7687 9255 7713
rect 9281 7687 9282 7713
rect 9254 7681 9282 7687
rect 9310 7938 9338 7943
rect 8862 7345 8890 7350
rect 9310 7321 9338 7910
rect 9366 7937 9394 7943
rect 9366 7911 9367 7937
rect 9393 7911 9394 7937
rect 9366 7713 9394 7911
rect 9366 7687 9367 7713
rect 9393 7687 9394 7713
rect 9366 7681 9394 7687
rect 9478 7714 9506 8134
rect 9478 7681 9506 7686
rect 9534 8162 9562 8167
rect 9534 7658 9562 8134
rect 9590 8049 9618 8302
rect 9814 8162 9842 8167
rect 9814 8115 9842 8134
rect 9926 8161 9954 8471
rect 9926 8135 9927 8161
rect 9953 8135 9954 8161
rect 9926 8129 9954 8135
rect 9982 8498 10010 8503
rect 9982 8106 10010 8470
rect 10150 8442 10178 9030
rect 10206 9025 10234 9030
rect 10598 9226 10626 9231
rect 10598 8946 10626 9198
rect 10598 8913 10626 8918
rect 10654 8722 10682 8727
rect 10598 8721 10682 8722
rect 10598 8695 10655 8721
rect 10681 8695 10682 8721
rect 10598 8694 10682 8695
rect 10598 8498 10626 8694
rect 10654 8689 10682 8694
rect 10766 8610 10794 9310
rect 10822 9170 10850 9175
rect 10822 8833 10850 9142
rect 10822 8807 10823 8833
rect 10849 8807 10850 8833
rect 10822 8801 10850 8807
rect 10710 8554 10738 8559
rect 10766 8554 10794 8582
rect 10710 8553 10794 8554
rect 10710 8527 10711 8553
rect 10737 8527 10794 8553
rect 10710 8526 10794 8527
rect 10710 8521 10738 8526
rect 10094 8441 10178 8442
rect 10094 8415 10151 8441
rect 10177 8415 10178 8441
rect 10094 8414 10178 8415
rect 10038 8386 10066 8391
rect 10038 8339 10066 8358
rect 10038 8106 10066 8111
rect 9982 8105 10066 8106
rect 9982 8079 10039 8105
rect 10065 8079 10066 8105
rect 9982 8078 10066 8079
rect 10038 8073 10066 8078
rect 9590 8023 9591 8049
rect 9617 8023 9618 8049
rect 9590 7994 9618 8023
rect 9590 7961 9618 7966
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9534 7625 9562 7630
rect 10094 7657 10122 8414
rect 10150 8409 10178 8414
rect 10430 8442 10458 8447
rect 10430 8395 10458 8414
rect 10598 8441 10626 8470
rect 10598 8415 10599 8441
rect 10625 8415 10626 8441
rect 10598 8330 10626 8415
rect 10878 8441 10906 9926
rect 11046 9921 11074 9926
rect 10990 9898 11018 9903
rect 10934 9870 10990 9898
rect 10934 9281 10962 9870
rect 10990 9865 11018 9870
rect 10990 9618 11018 9623
rect 10990 9337 11018 9590
rect 10990 9311 10991 9337
rect 11017 9311 11018 9337
rect 10990 9305 11018 9311
rect 10934 9255 10935 9281
rect 10961 9255 10962 9281
rect 10934 9249 10962 9255
rect 11270 9226 11298 11103
rect 11326 10850 11354 11662
rect 11382 11241 11410 11886
rect 11494 11858 11522 11863
rect 11494 11811 11522 11830
rect 11382 11215 11383 11241
rect 11409 11215 11410 11241
rect 11382 11209 11410 11215
rect 11550 11410 11578 11415
rect 11438 11129 11466 11135
rect 11438 11103 11439 11129
rect 11465 11103 11466 11129
rect 11438 10906 11466 11103
rect 11438 10873 11466 10878
rect 11326 9953 11354 10822
rect 11382 10737 11410 10743
rect 11382 10711 11383 10737
rect 11409 10711 11410 10737
rect 11382 10402 11410 10711
rect 11382 10355 11410 10374
rect 11550 10065 11578 11382
rect 11606 11130 11634 11135
rect 11606 11073 11634 11102
rect 11606 11047 11607 11073
rect 11633 11047 11634 11073
rect 11606 10570 11634 11047
rect 11718 11074 11746 11943
rect 11886 11969 11914 12334
rect 11886 11943 11887 11969
rect 11913 11943 11914 11969
rect 11886 11937 11914 11943
rect 11942 11858 11970 11863
rect 11942 11811 11970 11830
rect 11998 11857 12026 12390
rect 12334 12362 12362 12367
rect 12334 12305 12362 12334
rect 12334 12279 12335 12305
rect 12361 12279 12362 12305
rect 12334 12273 12362 12279
rect 11998 11831 11999 11857
rect 12025 11831 12026 11857
rect 11774 11074 11802 11079
rect 11718 11073 11802 11074
rect 11718 11047 11775 11073
rect 11801 11047 11802 11073
rect 11718 11046 11802 11047
rect 11662 10794 11690 10799
rect 11718 10794 11746 11046
rect 11774 11041 11802 11046
rect 11690 10766 11746 10794
rect 11662 10761 11690 10766
rect 11606 10542 11690 10570
rect 11550 10039 11551 10065
rect 11577 10039 11578 10065
rect 11326 9927 11327 9953
rect 11353 9927 11354 9953
rect 11326 9921 11354 9927
rect 11494 9954 11522 9959
rect 11326 9674 11354 9679
rect 11326 9627 11354 9646
rect 11494 9617 11522 9926
rect 11550 9898 11578 10039
rect 11662 9954 11690 10542
rect 11662 9921 11690 9926
rect 11718 10009 11746 10015
rect 11718 9983 11719 10009
rect 11745 9983 11746 10009
rect 11550 9865 11578 9870
rect 11494 9591 11495 9617
rect 11521 9591 11522 9617
rect 11494 9585 11522 9591
rect 11718 9674 11746 9983
rect 11718 9338 11746 9646
rect 11830 9617 11858 9623
rect 11830 9591 11831 9617
rect 11857 9591 11858 9617
rect 11718 9310 11802 9338
rect 11270 9193 11298 9198
rect 11662 9226 11690 9231
rect 10990 9114 11018 9119
rect 10990 9113 11074 9114
rect 10990 9087 10991 9113
rect 11017 9087 11074 9113
rect 10990 9086 11074 9087
rect 10990 9081 11018 9086
rect 10878 8415 10879 8441
rect 10905 8415 10906 8441
rect 10878 8409 10906 8415
rect 10598 8297 10626 8302
rect 10654 8385 10682 8391
rect 10654 8359 10655 8385
rect 10681 8359 10682 8385
rect 10654 8162 10682 8359
rect 10934 8386 10962 8391
rect 10934 8339 10962 8358
rect 10150 8134 10682 8162
rect 11046 8162 11074 9086
rect 11214 8722 11242 8727
rect 11158 8554 11186 8559
rect 11102 8526 11158 8554
rect 11102 8497 11130 8526
rect 11158 8521 11186 8526
rect 11102 8471 11103 8497
rect 11129 8471 11130 8497
rect 11102 8465 11130 8471
rect 11214 8497 11242 8694
rect 11662 8666 11690 9198
rect 11718 9225 11746 9231
rect 11718 9199 11719 9225
rect 11745 9199 11746 9225
rect 11718 9170 11746 9199
rect 11718 9137 11746 9142
rect 11774 8834 11802 9310
rect 11830 9170 11858 9591
rect 11886 9281 11914 9287
rect 11886 9255 11887 9281
rect 11913 9255 11914 9281
rect 11886 9226 11914 9255
rect 11886 9193 11914 9198
rect 11830 9137 11858 9142
rect 11886 8946 11914 8951
rect 11886 8899 11914 8918
rect 11886 8834 11914 8839
rect 11774 8833 11914 8834
rect 11774 8807 11887 8833
rect 11913 8807 11914 8833
rect 11774 8806 11914 8807
rect 11718 8778 11746 8783
rect 11718 8731 11746 8750
rect 11662 8638 11746 8666
rect 11550 8610 11578 8615
rect 11550 8553 11578 8582
rect 11550 8527 11551 8553
rect 11577 8527 11578 8553
rect 11550 8521 11578 8527
rect 11606 8554 11634 8559
rect 11606 8507 11634 8526
rect 11214 8471 11215 8497
rect 11241 8471 11242 8497
rect 11214 8442 11242 8471
rect 11662 8498 11690 8503
rect 11662 8451 11690 8470
rect 11214 8409 11242 8414
rect 11270 8441 11298 8447
rect 11270 8415 11271 8441
rect 11297 8415 11298 8441
rect 10150 8049 10178 8134
rect 11046 8129 11074 8134
rect 10150 8023 10151 8049
rect 10177 8023 10178 8049
rect 10150 8017 10178 8023
rect 10206 7938 10234 7943
rect 10206 7891 10234 7910
rect 10262 7938 10290 7943
rect 10262 7937 10346 7938
rect 10262 7911 10263 7937
rect 10289 7911 10346 7937
rect 10262 7910 10346 7911
rect 10262 7905 10290 7910
rect 10318 7713 10346 7910
rect 10318 7687 10319 7713
rect 10345 7687 10346 7713
rect 10318 7681 10346 7687
rect 10374 7714 10402 7719
rect 10374 7667 10402 7686
rect 11270 7713 11298 8415
rect 11326 8441 11354 8447
rect 11326 8415 11327 8441
rect 11353 8415 11354 8441
rect 11326 8162 11354 8415
rect 11326 7994 11354 8134
rect 11718 8161 11746 8638
rect 11774 8442 11802 8447
rect 11774 8441 11858 8442
rect 11774 8415 11775 8441
rect 11801 8415 11858 8441
rect 11774 8414 11858 8415
rect 11774 8409 11802 8414
rect 11718 8135 11719 8161
rect 11745 8135 11746 8161
rect 11718 8129 11746 8135
rect 11774 8330 11802 8335
rect 11774 8161 11802 8302
rect 11774 8135 11775 8161
rect 11801 8135 11802 8161
rect 11774 8129 11802 8135
rect 11830 8106 11858 8414
rect 11886 8441 11914 8806
rect 11998 8778 12026 11831
rect 12446 11857 12474 13454
rect 20118 13425 20146 13431
rect 20118 13399 20119 13425
rect 20145 13399 20146 13425
rect 13454 13202 13482 13207
rect 13454 13155 13482 13174
rect 12894 13146 12922 13151
rect 12894 13099 12922 13118
rect 13342 13146 13370 13151
rect 12782 13089 12810 13095
rect 12782 13063 12783 13089
rect 12809 13063 12810 13089
rect 12726 13034 12754 13039
rect 12614 13033 12754 13034
rect 12614 13007 12727 13033
rect 12753 13007 12754 13033
rect 12614 13006 12754 13007
rect 12614 12418 12642 13006
rect 12726 13001 12754 13006
rect 12782 12810 12810 13063
rect 13342 12810 13370 13118
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 20118 13146 20146 13399
rect 20118 13113 20146 13118
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 13454 12810 13482 12815
rect 13342 12809 13482 12810
rect 13342 12783 13455 12809
rect 13481 12783 13482 12809
rect 13342 12782 13482 12783
rect 12782 12777 12810 12782
rect 13454 12754 13482 12782
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 13454 12721 13482 12726
rect 18830 12754 18858 12759
rect 18830 12707 18858 12726
rect 13678 12642 13706 12647
rect 13678 12595 13706 12614
rect 13398 12586 13426 12591
rect 12614 12385 12642 12390
rect 12782 12418 12810 12423
rect 12782 12371 12810 12390
rect 12670 12362 12698 12367
rect 12670 12315 12698 12334
rect 12446 11831 12447 11857
rect 12473 11831 12474 11857
rect 12446 11802 12474 11831
rect 12446 11769 12474 11774
rect 13118 11690 13146 11695
rect 13118 11577 13146 11662
rect 13398 11690 13426 12558
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 18830 12194 18858 12199
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 18830 11969 18858 12166
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 18830 11943 18831 11969
rect 18857 11943 18858 11969
rect 18830 11937 18858 11943
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 13398 11657 13426 11662
rect 14798 11690 14826 11695
rect 14798 11643 14826 11662
rect 13118 11551 13119 11577
rect 13145 11551 13146 11577
rect 13118 10906 13146 11551
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 13510 11522 13538 11527
rect 13454 11521 13538 11522
rect 13454 11495 13511 11521
rect 13537 11495 13538 11521
rect 13454 11494 13538 11495
rect 13174 11242 13202 11247
rect 13174 11074 13202 11214
rect 13454 11241 13482 11494
rect 13510 11489 13538 11494
rect 13790 11522 13818 11527
rect 13454 11215 13455 11241
rect 13481 11215 13482 11241
rect 13454 11209 13482 11215
rect 13510 11186 13538 11191
rect 13734 11186 13762 11191
rect 13510 11185 13762 11186
rect 13510 11159 13511 11185
rect 13537 11159 13735 11185
rect 13761 11159 13762 11185
rect 13510 11158 13762 11159
rect 13510 11153 13538 11158
rect 13734 11153 13762 11158
rect 13790 11185 13818 11494
rect 14574 11522 14602 11527
rect 14574 11475 14602 11494
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 13790 11159 13791 11185
rect 13817 11159 13818 11185
rect 13790 11153 13818 11159
rect 14014 11186 14042 11191
rect 14014 11185 14210 11186
rect 14014 11159 14015 11185
rect 14041 11159 14210 11185
rect 14014 11158 14210 11159
rect 14014 11153 14042 11158
rect 13174 11027 13202 11046
rect 13398 11073 13426 11079
rect 13398 11047 13399 11073
rect 13425 11047 13426 11073
rect 13118 10873 13146 10878
rect 13342 10906 13370 10911
rect 12670 10850 12698 10855
rect 12670 10849 12754 10850
rect 12670 10823 12671 10849
rect 12697 10823 12754 10849
rect 12670 10822 12754 10823
rect 12670 10817 12698 10822
rect 12614 10793 12642 10799
rect 12614 10767 12615 10793
rect 12641 10767 12642 10793
rect 12614 10178 12642 10767
rect 12558 10150 12642 10178
rect 12670 10681 12698 10687
rect 12670 10655 12671 10681
rect 12697 10655 12698 10681
rect 12166 9954 12194 9959
rect 12166 9673 12194 9926
rect 12166 9647 12167 9673
rect 12193 9647 12194 9673
rect 12166 9641 12194 9647
rect 12558 9562 12586 10150
rect 12614 10066 12642 10071
rect 12670 10066 12698 10655
rect 12614 10065 12698 10066
rect 12614 10039 12615 10065
rect 12641 10039 12698 10065
rect 12614 10038 12698 10039
rect 12726 10066 12754 10822
rect 13342 10737 13370 10878
rect 13342 10711 13343 10737
rect 13369 10711 13370 10737
rect 12614 10033 12642 10038
rect 12726 10033 12754 10038
rect 13230 10066 13258 10071
rect 12782 10009 12810 10015
rect 12782 9983 12783 10009
rect 12809 9983 12810 10009
rect 12670 9954 12698 9959
rect 12670 9907 12698 9926
rect 12782 9730 12810 9983
rect 12838 10010 12866 10015
rect 12866 9982 12978 10010
rect 12838 9963 12866 9982
rect 12782 9697 12810 9702
rect 12334 9170 12362 9175
rect 12334 8834 12362 9142
rect 12334 8801 12362 8806
rect 11998 8745 12026 8750
rect 11886 8415 11887 8441
rect 11913 8415 11914 8441
rect 11886 8409 11914 8415
rect 11830 8078 12250 8106
rect 11326 7961 11354 7966
rect 11606 8049 11634 8055
rect 11606 8023 11607 8049
rect 11633 8023 11634 8049
rect 11270 7687 11271 7713
rect 11297 7687 11298 7713
rect 11270 7681 11298 7687
rect 10094 7631 10095 7657
rect 10121 7631 10122 7657
rect 10094 7625 10122 7631
rect 10206 7658 10234 7663
rect 10206 7611 10234 7630
rect 10934 7657 10962 7663
rect 10934 7631 10935 7657
rect 10961 7631 10962 7657
rect 10934 7574 10962 7631
rect 11606 7658 11634 8023
rect 11998 7993 12026 7999
rect 11998 7967 11999 7993
rect 12025 7967 12026 7993
rect 11774 7938 11802 7943
rect 11998 7938 12026 7967
rect 12110 7994 12138 7999
rect 12110 7947 12138 7966
rect 11774 7937 12026 7938
rect 11774 7911 11775 7937
rect 11801 7911 12026 7937
rect 11774 7910 12026 7911
rect 12166 7937 12194 7943
rect 12166 7911 12167 7937
rect 12193 7911 12194 7937
rect 11774 7905 11802 7910
rect 11606 7625 11634 7630
rect 11550 7602 11578 7607
rect 10486 7545 10514 7551
rect 10934 7546 11242 7574
rect 10486 7519 10487 7545
rect 10513 7519 10514 7545
rect 9310 7295 9311 7321
rect 9337 7295 9338 7321
rect 9310 7289 9338 7295
rect 9534 7322 9562 7327
rect 8918 7266 8946 7271
rect 8806 7265 8946 7266
rect 8806 7239 8919 7265
rect 8945 7239 8946 7265
rect 8806 7238 8946 7239
rect 8918 6985 8946 7238
rect 8918 6959 8919 6985
rect 8945 6959 8946 6985
rect 8918 6953 8946 6959
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 9534 2169 9562 7294
rect 10374 7322 10402 7327
rect 10486 7322 10514 7519
rect 10374 7321 10514 7322
rect 10374 7295 10375 7321
rect 10401 7295 10514 7321
rect 10374 7294 10514 7295
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10374 4214 10402 7294
rect 11214 7266 11242 7546
rect 11550 7266 11578 7574
rect 12166 7546 12194 7911
rect 12222 7574 12250 8078
rect 12558 8049 12586 9534
rect 12950 9225 12978 9982
rect 13230 9674 13258 10038
rect 13230 9627 13258 9646
rect 13342 9953 13370 10711
rect 13398 10738 13426 11047
rect 13678 11074 13706 11079
rect 13398 10705 13426 10710
rect 13566 10906 13594 10911
rect 13566 10793 13594 10878
rect 13566 10767 13567 10793
rect 13593 10767 13594 10793
rect 13566 10457 13594 10767
rect 13566 10431 13567 10457
rect 13593 10431 13594 10457
rect 13566 10425 13594 10431
rect 13622 10122 13650 10127
rect 13510 10066 13538 10071
rect 13510 10019 13538 10038
rect 13622 10065 13650 10094
rect 13622 10039 13623 10065
rect 13649 10039 13650 10065
rect 13622 10033 13650 10039
rect 13342 9927 13343 9953
rect 13369 9927 13370 9953
rect 13006 9338 13034 9343
rect 13006 9337 13258 9338
rect 13006 9311 13007 9337
rect 13033 9311 13258 9337
rect 13006 9310 13258 9311
rect 13006 9305 13034 9310
rect 12950 9199 12951 9225
rect 12977 9199 12978 9225
rect 12950 9193 12978 9199
rect 12838 9113 12866 9119
rect 12838 9087 12839 9113
rect 12865 9087 12866 9113
rect 12838 8946 12866 9087
rect 12838 8913 12866 8918
rect 13006 9113 13034 9119
rect 13006 9087 13007 9113
rect 13033 9087 13034 9113
rect 12558 8023 12559 8049
rect 12585 8023 12586 8049
rect 12558 8017 12586 8023
rect 12894 8834 12922 8839
rect 12278 7994 12306 7999
rect 12390 7994 12418 7999
rect 12278 7993 12418 7994
rect 12278 7967 12279 7993
rect 12305 7967 12391 7993
rect 12417 7967 12418 7993
rect 12278 7966 12418 7967
rect 12278 7961 12306 7966
rect 12390 7961 12418 7966
rect 12502 7938 12530 7943
rect 12502 7891 12530 7910
rect 12670 7657 12698 7663
rect 12670 7631 12671 7657
rect 12697 7631 12698 7657
rect 12334 7601 12362 7607
rect 12334 7575 12335 7601
rect 12361 7575 12362 7601
rect 12334 7574 12362 7575
rect 12222 7546 12362 7574
rect 12614 7602 12642 7607
rect 12670 7602 12698 7631
rect 12642 7574 12698 7602
rect 12894 7602 12922 8806
rect 13006 8386 13034 9087
rect 13230 8889 13258 9310
rect 13230 8863 13231 8889
rect 13257 8863 13258 8889
rect 13230 8857 13258 8863
rect 13286 9226 13314 9231
rect 13342 9226 13370 9927
rect 13678 9730 13706 11046
rect 13902 10738 13930 10743
rect 13734 10737 13930 10738
rect 13734 10711 13903 10737
rect 13929 10711 13930 10737
rect 13734 10710 13930 10711
rect 13734 10121 13762 10710
rect 13902 10705 13930 10710
rect 14182 10401 14210 11158
rect 18942 11185 18970 11191
rect 18942 11159 18943 11185
rect 18969 11159 18970 11185
rect 15302 10850 15330 10855
rect 15302 10803 15330 10822
rect 15190 10794 15218 10799
rect 14966 10766 15190 10794
rect 14966 10738 14994 10766
rect 15190 10747 15218 10766
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 14910 10737 14994 10738
rect 14910 10711 14967 10737
rect 14993 10711 14994 10737
rect 14910 10710 14994 10711
rect 14182 10375 14183 10401
rect 14209 10375 14210 10401
rect 13734 10095 13735 10121
rect 13761 10095 13762 10121
rect 13734 10089 13762 10095
rect 13846 10290 13874 10295
rect 13846 10009 13874 10262
rect 14182 10094 14210 10375
rect 14238 10402 14266 10407
rect 14238 10345 14266 10374
rect 14910 10402 14938 10710
rect 14966 10705 14994 10710
rect 18830 10626 18858 10631
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 14910 10355 14938 10374
rect 18830 10401 18858 10598
rect 18830 10375 18831 10401
rect 18857 10375 18858 10401
rect 18830 10369 18858 10375
rect 14238 10319 14239 10345
rect 14265 10319 14266 10345
rect 14238 10313 14266 10319
rect 15022 10346 15050 10351
rect 15022 10299 15050 10318
rect 18942 10346 18970 11159
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 20006 10794 20034 10799
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 20006 10458 20034 10463
rect 20006 10411 20034 10430
rect 18942 10313 18970 10318
rect 14350 10290 14378 10295
rect 14350 10243 14378 10262
rect 13846 9983 13847 10009
rect 13873 9983 13874 10009
rect 13846 9977 13874 9983
rect 13958 10066 14210 10094
rect 20006 10066 20034 10071
rect 13678 9702 13818 9730
rect 13286 9225 13370 9226
rect 13286 9199 13287 9225
rect 13313 9199 13370 9225
rect 13286 9198 13370 9199
rect 13398 9617 13426 9623
rect 13398 9591 13399 9617
rect 13425 9591 13426 9617
rect 13286 8834 13314 9198
rect 13398 8946 13426 9591
rect 13734 9618 13762 9623
rect 13790 9618 13818 9702
rect 13734 9617 13818 9618
rect 13734 9591 13735 9617
rect 13761 9591 13818 9617
rect 13734 9590 13818 9591
rect 13846 9618 13874 9623
rect 13566 9562 13594 9567
rect 13734 9562 13762 9590
rect 13846 9571 13874 9590
rect 13566 9561 13706 9562
rect 13566 9535 13567 9561
rect 13593 9535 13706 9561
rect 13566 9534 13706 9535
rect 13566 9529 13594 9534
rect 13510 9505 13538 9511
rect 13510 9479 13511 9505
rect 13537 9479 13538 9505
rect 13510 9338 13538 9479
rect 13678 9450 13706 9534
rect 13734 9529 13762 9534
rect 13790 9505 13818 9511
rect 13790 9479 13791 9505
rect 13817 9479 13818 9505
rect 13790 9450 13818 9479
rect 13678 9422 13818 9450
rect 13958 9505 13986 10066
rect 18830 10009 18858 10015
rect 18830 9983 18831 10009
rect 18857 9983 18858 10009
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 18830 9730 18858 9983
rect 20006 9953 20034 10038
rect 20006 9927 20007 9953
rect 20033 9927 20034 9953
rect 20006 9921 20034 9927
rect 18830 9697 18858 9702
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 14686 9618 14714 9623
rect 14238 9562 14266 9567
rect 14238 9515 14266 9534
rect 13958 9479 13959 9505
rect 13985 9479 13986 9505
rect 13510 9310 13650 9338
rect 13622 9281 13650 9310
rect 13622 9255 13623 9281
rect 13649 9255 13650 9281
rect 13622 9249 13650 9255
rect 13958 9226 13986 9479
rect 13958 9193 13986 9198
rect 14686 9169 14714 9590
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 14686 9143 14687 9169
rect 14713 9143 14714 9169
rect 14686 9137 14714 9143
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 13398 8913 13426 8918
rect 13286 8801 13314 8806
rect 13566 8890 13594 8895
rect 13398 8778 13426 8783
rect 13398 8497 13426 8750
rect 13398 8471 13399 8497
rect 13425 8471 13426 8497
rect 13398 8465 13426 8471
rect 13566 8441 13594 8862
rect 14294 8890 14322 8895
rect 14294 8843 14322 8862
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 14630 8834 14658 8839
rect 14630 8787 14658 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 13566 8415 13567 8441
rect 13593 8415 13594 8441
rect 13566 8409 13594 8415
rect 13006 8353 13034 8358
rect 13454 8386 13482 8391
rect 13454 8339 13482 8358
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 12614 7569 12642 7574
rect 12894 7569 12922 7574
rect 13006 7938 13034 7943
rect 11942 7518 12194 7546
rect 11942 7321 11970 7518
rect 11942 7295 11943 7321
rect 11969 7295 11970 7321
rect 11942 7289 11970 7295
rect 11214 7265 11578 7266
rect 11214 7239 11551 7265
rect 11577 7239 11578 7265
rect 11214 7238 11578 7239
rect 11550 7233 11578 7238
rect 12334 4214 12362 7546
rect 13006 7321 13034 7910
rect 13006 7295 13007 7321
rect 13033 7295 13034 7321
rect 13006 4214 13034 7295
rect 13286 7602 13314 7607
rect 13286 7321 13314 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13286 7295 13287 7321
rect 13313 7295 13314 7321
rect 13286 7289 13314 7295
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 10374 4186 10570 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9534 2143 9535 2169
rect 9561 2143 9562 2169
rect 9534 2137 9562 2143
rect 9422 2058 9450 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 9422 400 9450 2030
rect 10038 2058 10066 2063
rect 10038 2011 10066 2030
rect 10430 1834 10458 1839
rect 10094 1665 10122 1671
rect 10094 1639 10095 1665
rect 10121 1639 10122 1665
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10094 400 10122 1639
rect 10430 400 10458 1806
rect 10542 1777 10570 4186
rect 12278 4186 12362 4214
rect 12614 4186 13034 4214
rect 11046 1834 11074 1839
rect 11046 1787 11074 1806
rect 11438 1834 11466 1839
rect 10542 1751 10543 1777
rect 10569 1751 10570 1777
rect 10542 1745 10570 1751
rect 11438 400 11466 1806
rect 12278 1777 12306 4186
rect 12614 2169 12642 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12446 2058 12474 2063
rect 12446 400 12474 2030
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 9408 0 9464 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 11424 0 11480 400
rect 12432 0 12488 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 8750 14238 8778 14266
rect 2086 13790 2114 13818
rect 966 13118 994 13146
rect 966 12782 994 12810
rect 966 11774 994 11802
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2142 13454 2170 13482
rect 5782 13454 5810 13482
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 5726 13118 5754 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 7462 13481 7490 13482
rect 7462 13455 7463 13481
rect 7463 13455 7489 13481
rect 7489 13455 7490 13481
rect 7462 13454 7490 13455
rect 6846 13145 6874 13146
rect 6846 13119 6847 13145
rect 6847 13119 6873 13145
rect 6873 13119 6874 13145
rect 6846 13118 6874 13119
rect 5726 12670 5754 12698
rect 6902 12726 6930 12754
rect 7630 13398 7658 13426
rect 7798 13145 7826 13146
rect 7798 13119 7799 13145
rect 7799 13119 7825 13145
rect 7825 13119 7826 13145
rect 7798 13118 7826 13119
rect 7742 13062 7770 13090
rect 7462 13033 7490 13034
rect 7462 13007 7463 13033
rect 7463 13007 7489 13033
rect 7489 13007 7490 13033
rect 7462 13006 7490 13007
rect 7350 12726 7378 12754
rect 7406 12782 7434 12810
rect 7350 12641 7378 12642
rect 7350 12615 7351 12641
rect 7351 12615 7377 12641
rect 7377 12615 7378 12641
rect 7350 12614 7378 12615
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 6510 11942 6538 11970
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 4942 11494 4970 11522
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6286 11521 6314 11522
rect 6286 11495 6287 11521
rect 6287 11495 6313 11521
rect 6313 11495 6314 11521
rect 6286 11494 6314 11495
rect 2086 11046 2114 11074
rect 5334 10878 5362 10906
rect 6342 10934 6370 10962
rect 6006 10822 6034 10850
rect 6510 11102 6538 11130
rect 7014 11718 7042 11746
rect 7014 10990 7042 11018
rect 6790 10934 6818 10962
rect 6398 10766 6426 10794
rect 5670 10737 5698 10738
rect 5670 10711 5671 10737
rect 5671 10711 5697 10737
rect 5697 10711 5698 10737
rect 5670 10710 5698 10711
rect 6734 10654 6762 10682
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6958 10793 6986 10794
rect 6958 10767 6959 10793
rect 6959 10767 6985 10793
rect 6985 10767 6986 10793
rect 6958 10766 6986 10767
rect 7854 12697 7882 12698
rect 7854 12671 7855 12697
rect 7855 12671 7881 12697
rect 7881 12671 7882 12697
rect 7854 12670 7882 12671
rect 8134 13230 8162 13258
rect 8694 13566 8722 13594
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12110 19110 12138 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9758 18718 9786 18746
rect 10374 18745 10402 18746
rect 10374 18719 10375 18745
rect 10375 18719 10401 18745
rect 10401 18719 10402 18745
rect 10374 18718 10402 18719
rect 9366 14265 9394 14266
rect 9366 14239 9367 14265
rect 9367 14239 9393 14265
rect 9393 14239 9394 14265
rect 9366 14238 9394 14239
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9478 14265 9506 14266
rect 9478 14239 9479 14265
rect 9479 14239 9505 14265
rect 9505 14239 9506 14265
rect 9478 14238 9506 14239
rect 9422 13622 9450 13650
rect 8862 13257 8890 13258
rect 8862 13231 8863 13257
rect 8863 13231 8889 13257
rect 8889 13231 8890 13257
rect 8862 13230 8890 13231
rect 10150 14238 10178 14266
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9814 13902 9842 13930
rect 9758 13593 9786 13594
rect 9758 13567 9759 13593
rect 9759 13567 9785 13593
rect 9785 13567 9786 13593
rect 9758 13566 9786 13567
rect 7910 12614 7938 12642
rect 7462 11718 7490 11746
rect 7574 11633 7602 11634
rect 7574 11607 7575 11633
rect 7575 11607 7601 11633
rect 7601 11607 7602 11633
rect 7574 11606 7602 11607
rect 7406 10934 7434 10962
rect 7518 11494 7546 11522
rect 7350 10905 7378 10906
rect 7350 10879 7351 10905
rect 7351 10879 7377 10905
rect 7377 10879 7378 10905
rect 7350 10878 7378 10879
rect 7182 10849 7210 10850
rect 7182 10823 7183 10849
rect 7183 10823 7209 10849
rect 7209 10823 7210 10849
rect 7182 10822 7210 10823
rect 7294 10793 7322 10794
rect 7294 10767 7295 10793
rect 7295 10767 7321 10793
rect 7321 10767 7322 10793
rect 7294 10766 7322 10767
rect 6846 10457 6874 10458
rect 6846 10431 6847 10457
rect 6847 10431 6873 10457
rect 6873 10431 6874 10457
rect 6846 10430 6874 10431
rect 4998 9982 5026 10010
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 4998 9673 5026 9674
rect 4998 9647 4999 9673
rect 4999 9647 5025 9673
rect 5025 9647 5026 9673
rect 4998 9646 5026 9647
rect 2142 9617 2170 9618
rect 2142 9591 2143 9617
rect 2143 9591 2169 9617
rect 2169 9591 2170 9617
rect 2142 9590 2170 9591
rect 6454 9617 6482 9618
rect 6454 9591 6455 9617
rect 6455 9591 6481 9617
rect 6481 9591 6482 9617
rect 6454 9590 6482 9591
rect 7126 10009 7154 10010
rect 7126 9983 7127 10009
rect 7127 9983 7153 10009
rect 7153 9983 7154 10009
rect 7126 9982 7154 9983
rect 6790 9590 6818 9618
rect 966 9422 994 9450
rect 6062 9310 6090 9338
rect 6734 9534 6762 9562
rect 6678 9086 6706 9114
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 5838 8497 5866 8498
rect 5838 8471 5839 8497
rect 5839 8471 5865 8497
rect 5865 8471 5866 8497
rect 5838 8470 5866 8471
rect 5502 8441 5530 8442
rect 5502 8415 5503 8441
rect 5503 8415 5529 8441
rect 5529 8415 5530 8441
rect 5502 8414 5530 8415
rect 6342 8358 6370 8386
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 7126 9534 7154 9562
rect 6958 9225 6986 9226
rect 6958 9199 6959 9225
rect 6959 9199 6985 9225
rect 6985 9199 6986 9225
rect 6958 9198 6986 9199
rect 6902 9169 6930 9170
rect 6902 9143 6903 9169
rect 6903 9143 6929 9169
rect 6929 9143 6930 9169
rect 6902 9142 6930 9143
rect 7126 9337 7154 9338
rect 7126 9311 7127 9337
rect 7127 9311 7153 9337
rect 7153 9311 7154 9337
rect 7126 9310 7154 9311
rect 7406 10206 7434 10234
rect 7462 10150 7490 10178
rect 7574 10793 7602 10794
rect 7574 10767 7575 10793
rect 7575 10767 7601 10793
rect 7601 10767 7602 10793
rect 7574 10766 7602 10767
rect 7406 9870 7434 9898
rect 7238 9617 7266 9618
rect 7238 9591 7239 9617
rect 7239 9591 7265 9617
rect 7265 9591 7266 9617
rect 7238 9590 7266 9591
rect 7350 9478 7378 9506
rect 7182 9030 7210 9058
rect 7238 9086 7266 9114
rect 7910 11942 7938 11970
rect 8134 12334 8162 12362
rect 8078 11857 8106 11858
rect 8078 11831 8079 11857
rect 8079 11831 8105 11857
rect 8105 11831 8106 11857
rect 8078 11830 8106 11831
rect 8190 12782 8218 12810
rect 8806 13062 8834 13090
rect 9646 13145 9674 13146
rect 9646 13119 9647 13145
rect 9647 13119 9673 13145
rect 9673 13119 9674 13145
rect 9646 13118 9674 13119
rect 10654 13929 10682 13930
rect 10654 13903 10655 13929
rect 10655 13903 10681 13929
rect 10681 13903 10682 13929
rect 10654 13902 10682 13903
rect 10262 13678 10290 13706
rect 10150 13398 10178 13426
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9254 12614 9282 12642
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10374 13622 10402 13650
rect 11718 13846 11746 13874
rect 11438 13678 11466 13706
rect 11270 13622 11298 13650
rect 11158 13566 11186 13594
rect 10654 13454 10682 13482
rect 10878 13454 10906 13482
rect 9590 12417 9618 12418
rect 9590 12391 9591 12417
rect 9591 12391 9617 12417
rect 9617 12391 9618 12417
rect 9590 12390 9618 12391
rect 8470 11830 8498 11858
rect 8190 11718 8218 11746
rect 8694 11718 8722 11746
rect 8190 11633 8218 11634
rect 8190 11607 8191 11633
rect 8191 11607 8217 11633
rect 8217 11607 8218 11633
rect 8190 11606 8218 11607
rect 7798 11158 7826 11186
rect 7910 10934 7938 10962
rect 8078 11158 8106 11186
rect 8078 10934 8106 10962
rect 7686 10737 7714 10738
rect 7686 10711 7687 10737
rect 7687 10711 7713 10737
rect 7713 10711 7714 10737
rect 7686 10710 7714 10711
rect 7742 10457 7770 10458
rect 7742 10431 7743 10457
rect 7743 10431 7769 10457
rect 7769 10431 7770 10457
rect 7742 10430 7770 10431
rect 7462 9646 7490 9674
rect 7630 9617 7658 9618
rect 7630 9591 7631 9617
rect 7631 9591 7657 9617
rect 7657 9591 7658 9617
rect 7630 9590 7658 9591
rect 7742 9561 7770 9562
rect 7742 9535 7743 9561
rect 7743 9535 7769 9561
rect 7769 9535 7770 9561
rect 7742 9534 7770 9535
rect 7518 9281 7546 9282
rect 7518 9255 7519 9281
rect 7519 9255 7545 9281
rect 7545 9255 7546 9281
rect 7518 9254 7546 9255
rect 7462 9198 7490 9226
rect 7910 10710 7938 10738
rect 8022 10766 8050 10794
rect 8414 11577 8442 11578
rect 8414 11551 8415 11577
rect 8415 11551 8441 11577
rect 8441 11551 8442 11577
rect 8414 11550 8442 11551
rect 8694 11241 8722 11242
rect 8694 11215 8695 11241
rect 8695 11215 8721 11241
rect 8721 11215 8722 11241
rect 8694 11214 8722 11215
rect 8190 11129 8218 11130
rect 8190 11103 8191 11129
rect 8191 11103 8217 11129
rect 8217 11103 8218 11129
rect 8190 11102 8218 11103
rect 8246 10934 8274 10962
rect 8078 10206 8106 10234
rect 8190 10094 8218 10122
rect 7966 10038 7994 10066
rect 8302 10793 8330 10794
rect 8302 10767 8303 10793
rect 8303 10767 8329 10793
rect 8329 10767 8330 10793
rect 8302 10766 8330 10767
rect 7966 9590 7994 9618
rect 10206 12361 10234 12362
rect 10206 12335 10207 12361
rect 10207 12335 10233 12361
rect 10233 12335 10234 12361
rect 10206 12334 10234 12335
rect 8862 11577 8890 11578
rect 8862 11551 8863 11577
rect 8863 11551 8889 11577
rect 8889 11551 8890 11577
rect 8862 11550 8890 11551
rect 8750 11158 8778 11186
rect 8694 10766 8722 10794
rect 8470 10654 8498 10682
rect 8862 10654 8890 10682
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10374 11718 10402 11746
rect 9254 11550 9282 11578
rect 10038 11606 10066 11634
rect 9590 11521 9618 11522
rect 9590 11495 9591 11521
rect 9591 11495 9617 11521
rect 9617 11495 9618 11521
rect 9590 11494 9618 11495
rect 9310 11158 9338 11186
rect 9030 11102 9058 11130
rect 9086 11073 9114 11074
rect 9086 11047 9087 11073
rect 9087 11047 9113 11073
rect 9113 11047 9114 11073
rect 9086 11046 9114 11047
rect 9422 11129 9450 11130
rect 9422 11103 9423 11129
rect 9423 11103 9449 11129
rect 9449 11103 9450 11129
rect 9422 11102 9450 11103
rect 9198 10793 9226 10794
rect 9198 10767 9199 10793
rect 9199 10767 9225 10793
rect 9225 10767 9226 10793
rect 9198 10766 9226 10767
rect 6958 8470 6986 8498
rect 8414 10038 8442 10066
rect 8526 10206 8554 10234
rect 8134 9225 8162 9226
rect 8134 9199 8135 9225
rect 8135 9199 8161 9225
rect 8161 9199 8162 9225
rect 8134 9198 8162 9199
rect 8078 9086 8106 9114
rect 7966 8918 7994 8946
rect 7854 8694 7882 8722
rect 6790 8358 6818 8386
rect 6902 8414 6930 8442
rect 7350 8441 7378 8442
rect 7350 8415 7351 8441
rect 7351 8415 7377 8441
rect 7377 8415 7378 8441
rect 7350 8414 7378 8415
rect 7574 8414 7602 8442
rect 7630 8358 7658 8386
rect 8302 9534 8330 9562
rect 8358 10009 8386 10010
rect 8358 9983 8359 10009
rect 8359 9983 8385 10009
rect 8385 9983 8386 10009
rect 8358 9982 8386 9983
rect 8190 9086 8218 9114
rect 8246 9142 8274 9170
rect 8862 9729 8890 9730
rect 8862 9703 8863 9729
rect 8863 9703 8889 9729
rect 8889 9703 8890 9729
rect 8862 9702 8890 9703
rect 8974 9953 9002 9954
rect 8974 9927 8975 9953
rect 8975 9927 9001 9953
rect 9001 9927 9002 9953
rect 8974 9926 9002 9927
rect 8414 9198 8442 9226
rect 8246 8806 8274 8834
rect 8582 8833 8610 8834
rect 8582 8807 8583 8833
rect 8583 8807 8609 8833
rect 8609 8807 8610 8833
rect 8582 8806 8610 8807
rect 8918 9254 8946 9282
rect 8974 9225 9002 9226
rect 8974 9199 8975 9225
rect 8975 9199 9001 9225
rect 9001 9199 9002 9225
rect 8974 9198 9002 9199
rect 8806 8526 8834 8554
rect 7798 8414 7826 8442
rect 9254 10737 9282 10738
rect 9254 10711 9255 10737
rect 9255 10711 9281 10737
rect 9281 10711 9282 10737
rect 9254 10710 9282 10711
rect 9534 11046 9562 11074
rect 9590 10990 9618 11018
rect 9142 10318 9170 10346
rect 10318 11633 10346 11634
rect 10318 11607 10319 11633
rect 10319 11607 10345 11633
rect 10345 11607 10346 11633
rect 10318 11606 10346 11607
rect 10094 11550 10122 11578
rect 10094 11185 10122 11186
rect 10094 11159 10095 11185
rect 10095 11159 10121 11185
rect 10121 11159 10122 11185
rect 10094 11158 10122 11159
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9086 9617 9114 9618
rect 9086 9591 9087 9617
rect 9087 9591 9113 9617
rect 9113 9591 9114 9617
rect 9086 9590 9114 9591
rect 9198 9590 9226 9618
rect 9254 10206 9282 10234
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10038 10121 10066 10122
rect 10038 10095 10039 10121
rect 10039 10095 10065 10121
rect 10065 10095 10066 10121
rect 10038 10094 10066 10095
rect 9590 10065 9618 10066
rect 9590 10039 9591 10065
rect 9591 10039 9617 10065
rect 9617 10039 9618 10065
rect 9590 10038 9618 10039
rect 9366 9982 9394 10010
rect 9534 9926 9562 9954
rect 9310 8553 9338 8554
rect 9310 8527 9311 8553
rect 9311 8527 9337 8553
rect 9337 8527 9338 8553
rect 9310 8526 9338 8527
rect 9030 8414 9058 8442
rect 9254 8470 9282 8498
rect 7742 8161 7770 8162
rect 7742 8135 7743 8161
rect 7743 8135 7769 8161
rect 7769 8135 7770 8161
rect 7742 8134 7770 8135
rect 6678 7910 6706 7938
rect 6342 7574 6370 7602
rect 7686 7937 7714 7938
rect 7686 7911 7687 7937
rect 7687 7911 7713 7937
rect 7713 7911 7714 7937
rect 7686 7910 7714 7911
rect 7686 7686 7714 7714
rect 7014 7574 7042 7602
rect 7350 7574 7378 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8694 8134 8722 8162
rect 8806 7993 8834 7994
rect 8806 7967 8807 7993
rect 8807 7967 8833 7993
rect 8833 7967 8834 7993
rect 8806 7966 8834 7967
rect 7966 7601 7994 7602
rect 7966 7575 7967 7601
rect 7967 7575 7993 7601
rect 7993 7575 7994 7601
rect 7966 7574 7994 7575
rect 8750 7601 8778 7602
rect 8750 7575 8751 7601
rect 8751 7575 8777 7601
rect 8777 7575 8778 7601
rect 8750 7574 8778 7575
rect 8750 7321 8778 7322
rect 8750 7295 8751 7321
rect 8751 7295 8777 7321
rect 8777 7295 8778 7321
rect 8750 7294 8778 7295
rect 9142 7713 9170 7714
rect 9142 7687 9143 7713
rect 9143 7687 9169 7713
rect 9169 7687 9170 7713
rect 9142 7686 9170 7687
rect 9422 9534 9450 9562
rect 9814 10065 9842 10066
rect 9814 10039 9815 10065
rect 9815 10039 9841 10065
rect 9841 10039 9842 10065
rect 9814 10038 9842 10039
rect 9982 9982 10010 10010
rect 9758 9478 9786 9506
rect 10038 9505 10066 9506
rect 10038 9479 10039 9505
rect 10039 9479 10065 9505
rect 10065 9479 10066 9505
rect 10038 9478 10066 9479
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9814 9198 9842 9226
rect 11102 13398 11130 13426
rect 11662 13593 11690 13594
rect 11662 13567 11663 13593
rect 11663 13567 11689 13593
rect 11689 13567 11690 13593
rect 11662 13566 11690 13567
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 12110 13873 12138 13874
rect 12110 13847 12111 13873
rect 12111 13847 12137 13873
rect 12137 13847 12138 13873
rect 12110 13846 12138 13847
rect 12054 13454 12082 13482
rect 11550 13398 11578 13426
rect 11494 12782 11522 12810
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12390 13454 12418 13482
rect 11606 12697 11634 12698
rect 11606 12671 11607 12697
rect 11607 12671 11633 12697
rect 11633 12671 11634 12697
rect 11606 12670 11634 12671
rect 12390 12697 12418 12698
rect 12390 12671 12391 12697
rect 12391 12671 12417 12697
rect 12417 12671 12418 12697
rect 12390 12670 12418 12671
rect 11550 12641 11578 12642
rect 11550 12615 11551 12641
rect 11551 12615 11577 12641
rect 11577 12615 11578 12641
rect 11550 12614 11578 12615
rect 10654 11942 10682 11970
rect 10766 11718 10794 11746
rect 10822 11774 10850 11802
rect 10654 11577 10682 11578
rect 10654 11551 10655 11577
rect 10655 11551 10681 11577
rect 10681 11551 10682 11577
rect 10654 11550 10682 11551
rect 10766 11382 10794 11410
rect 10374 10934 10402 10962
rect 10206 10542 10234 10570
rect 10766 10934 10794 10962
rect 10766 10318 10794 10346
rect 10654 10262 10682 10290
rect 10262 10009 10290 10010
rect 10262 9983 10263 10009
rect 10263 9983 10289 10009
rect 10289 9983 10290 10009
rect 10262 9982 10290 9983
rect 10878 11185 10906 11186
rect 10878 11159 10879 11185
rect 10879 11159 10905 11185
rect 10905 11159 10906 11185
rect 10878 11158 10906 11159
rect 10934 10878 10962 10906
rect 10934 10542 10962 10570
rect 10878 10038 10906 10066
rect 11158 11969 11186 11970
rect 11158 11943 11159 11969
rect 11159 11943 11185 11969
rect 11185 11943 11186 11969
rect 11158 11942 11186 11943
rect 11270 12110 11298 12138
rect 11550 12110 11578 12138
rect 11998 12390 12026 12418
rect 11886 12334 11914 12362
rect 11270 11774 11298 11802
rect 11158 10934 11186 10962
rect 11102 10094 11130 10122
rect 11214 9982 11242 10010
rect 10654 9617 10682 9618
rect 10654 9591 10655 9617
rect 10655 9591 10681 9617
rect 10681 9591 10682 9617
rect 10654 9590 10682 9591
rect 10822 9561 10850 9562
rect 10822 9535 10823 9561
rect 10823 9535 10849 9561
rect 10849 9535 10850 9561
rect 10822 9534 10850 9535
rect 10766 9337 10794 9338
rect 10766 9311 10767 9337
rect 10767 9311 10793 9337
rect 10793 9311 10794 9337
rect 10766 9310 10794 9311
rect 10094 9142 10122 9170
rect 10206 9030 10234 9058
rect 9702 8806 9730 8834
rect 9366 8134 9394 8162
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9926 8526 9954 8554
rect 9814 8497 9842 8498
rect 9814 8471 9815 8497
rect 9815 8471 9841 8497
rect 9841 8471 9842 8497
rect 9814 8470 9842 8471
rect 9590 8302 9618 8330
rect 9310 7910 9338 7938
rect 8862 7350 8890 7378
rect 9478 7686 9506 7714
rect 9534 8161 9562 8162
rect 9534 8135 9535 8161
rect 9535 8135 9561 8161
rect 9561 8135 9562 8161
rect 9534 8134 9562 8135
rect 9814 8161 9842 8162
rect 9814 8135 9815 8161
rect 9815 8135 9841 8161
rect 9841 8135 9842 8161
rect 9814 8134 9842 8135
rect 9982 8470 10010 8498
rect 10598 9225 10626 9226
rect 10598 9199 10599 9225
rect 10599 9199 10625 9225
rect 10625 9199 10626 9225
rect 10598 9198 10626 9199
rect 10598 8918 10626 8946
rect 10822 9142 10850 9170
rect 10766 8582 10794 8610
rect 10598 8470 10626 8498
rect 10038 8385 10066 8386
rect 10038 8359 10039 8385
rect 10039 8359 10065 8385
rect 10065 8359 10066 8385
rect 10038 8358 10066 8359
rect 9590 7966 9618 7994
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9534 7630 9562 7658
rect 10430 8441 10458 8442
rect 10430 8415 10431 8441
rect 10431 8415 10457 8441
rect 10457 8415 10458 8441
rect 10430 8414 10458 8415
rect 11046 9926 11074 9954
rect 10990 9870 11018 9898
rect 10990 9590 11018 9618
rect 11494 11857 11522 11858
rect 11494 11831 11495 11857
rect 11495 11831 11521 11857
rect 11521 11831 11522 11857
rect 11494 11830 11522 11831
rect 11550 11382 11578 11410
rect 11438 10878 11466 10906
rect 11326 10822 11354 10850
rect 11382 10401 11410 10402
rect 11382 10375 11383 10401
rect 11383 10375 11409 10401
rect 11409 10375 11410 10401
rect 11382 10374 11410 10375
rect 11606 11102 11634 11130
rect 11942 11857 11970 11858
rect 11942 11831 11943 11857
rect 11943 11831 11969 11857
rect 11969 11831 11970 11857
rect 11942 11830 11970 11831
rect 12334 12334 12362 12362
rect 11662 10766 11690 10794
rect 11494 9926 11522 9954
rect 11326 9673 11354 9674
rect 11326 9647 11327 9673
rect 11327 9647 11353 9673
rect 11353 9647 11354 9673
rect 11326 9646 11354 9647
rect 11662 9926 11690 9954
rect 11550 9870 11578 9898
rect 11718 9646 11746 9674
rect 11270 9198 11298 9226
rect 11662 9198 11690 9226
rect 10598 8302 10626 8330
rect 10934 8385 10962 8386
rect 10934 8359 10935 8385
rect 10935 8359 10961 8385
rect 10961 8359 10962 8385
rect 10934 8358 10962 8359
rect 11214 8694 11242 8722
rect 11158 8526 11186 8554
rect 11718 9142 11746 9170
rect 11886 9198 11914 9226
rect 11830 9142 11858 9170
rect 11886 8945 11914 8946
rect 11886 8919 11887 8945
rect 11887 8919 11913 8945
rect 11913 8919 11914 8945
rect 11886 8918 11914 8919
rect 11718 8777 11746 8778
rect 11718 8751 11719 8777
rect 11719 8751 11745 8777
rect 11745 8751 11746 8777
rect 11718 8750 11746 8751
rect 11550 8582 11578 8610
rect 11606 8553 11634 8554
rect 11606 8527 11607 8553
rect 11607 8527 11633 8553
rect 11633 8527 11634 8553
rect 11606 8526 11634 8527
rect 11662 8497 11690 8498
rect 11662 8471 11663 8497
rect 11663 8471 11689 8497
rect 11689 8471 11690 8497
rect 11662 8470 11690 8471
rect 11214 8414 11242 8442
rect 11046 8134 11074 8162
rect 10206 7937 10234 7938
rect 10206 7911 10207 7937
rect 10207 7911 10233 7937
rect 10233 7911 10234 7937
rect 10206 7910 10234 7911
rect 10374 7713 10402 7714
rect 10374 7687 10375 7713
rect 10375 7687 10401 7713
rect 10401 7687 10402 7713
rect 10374 7686 10402 7687
rect 11326 8134 11354 8162
rect 11774 8302 11802 8330
rect 13454 13201 13482 13202
rect 13454 13175 13455 13201
rect 13455 13175 13481 13201
rect 13481 13175 13482 13201
rect 13454 13174 13482 13175
rect 12894 13145 12922 13146
rect 12894 13119 12895 13145
rect 12895 13119 12921 13145
rect 12921 13119 12922 13145
rect 12894 13118 12922 13119
rect 13342 13145 13370 13146
rect 13342 13119 13343 13145
rect 13343 13119 13369 13145
rect 13369 13119 13370 13145
rect 13342 13118 13370 13119
rect 12782 12782 12810 12810
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 20118 13118 20146 13146
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 19950 12782 19978 12810
rect 13454 12726 13482 12754
rect 18830 12753 18858 12754
rect 18830 12727 18831 12753
rect 18831 12727 18857 12753
rect 18857 12727 18858 12753
rect 18830 12726 18858 12727
rect 13678 12641 13706 12642
rect 13678 12615 13679 12641
rect 13679 12615 13705 12641
rect 13705 12615 13706 12641
rect 13678 12614 13706 12615
rect 13398 12558 13426 12586
rect 12614 12390 12642 12418
rect 12782 12417 12810 12418
rect 12782 12391 12783 12417
rect 12783 12391 12809 12417
rect 12809 12391 12810 12417
rect 12782 12390 12810 12391
rect 12670 12361 12698 12362
rect 12670 12335 12671 12361
rect 12671 12335 12697 12361
rect 12697 12335 12698 12361
rect 12670 12334 12698 12335
rect 12446 11774 12474 11802
rect 13118 11662 13146 11690
rect 20006 12446 20034 12474
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 18830 12166 18858 12194
rect 20006 12110 20034 12138
rect 20006 11774 20034 11802
rect 13398 11662 13426 11690
rect 14798 11689 14826 11690
rect 14798 11663 14799 11689
rect 14799 11663 14825 11689
rect 14825 11663 14826 11689
rect 14798 11662 14826 11663
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 13174 11214 13202 11242
rect 13790 11494 13818 11522
rect 14574 11521 14602 11522
rect 14574 11495 14575 11521
rect 14575 11495 14601 11521
rect 14601 11495 14602 11521
rect 14574 11494 14602 11495
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 13174 11073 13202 11074
rect 13174 11047 13175 11073
rect 13175 11047 13201 11073
rect 13201 11047 13202 11073
rect 13174 11046 13202 11047
rect 13118 10878 13146 10906
rect 13342 10878 13370 10906
rect 12166 9926 12194 9954
rect 12726 10038 12754 10066
rect 13230 10038 13258 10066
rect 12670 9953 12698 9954
rect 12670 9927 12671 9953
rect 12671 9927 12697 9953
rect 12697 9927 12698 9953
rect 12670 9926 12698 9927
rect 12838 10009 12866 10010
rect 12838 9983 12839 10009
rect 12839 9983 12865 10009
rect 12865 9983 12866 10009
rect 12838 9982 12866 9983
rect 12782 9702 12810 9730
rect 12558 9534 12586 9562
rect 12334 9169 12362 9170
rect 12334 9143 12335 9169
rect 12335 9143 12361 9169
rect 12361 9143 12362 9169
rect 12334 9142 12362 9143
rect 12334 8806 12362 8834
rect 11998 8750 12026 8778
rect 11326 7966 11354 7994
rect 10206 7657 10234 7658
rect 10206 7631 10207 7657
rect 10207 7631 10233 7657
rect 10233 7631 10234 7657
rect 10206 7630 10234 7631
rect 12110 7993 12138 7994
rect 12110 7967 12111 7993
rect 12111 7967 12137 7993
rect 12137 7967 12138 7993
rect 12110 7966 12138 7967
rect 11606 7630 11634 7658
rect 11550 7574 11578 7602
rect 9534 7294 9562 7322
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 13230 9673 13258 9674
rect 13230 9647 13231 9673
rect 13231 9647 13257 9673
rect 13257 9647 13258 9673
rect 13230 9646 13258 9647
rect 13678 11073 13706 11074
rect 13678 11047 13679 11073
rect 13679 11047 13705 11073
rect 13705 11047 13706 11073
rect 13678 11046 13706 11047
rect 13398 10710 13426 10738
rect 13566 10878 13594 10906
rect 13622 10094 13650 10122
rect 13510 10065 13538 10066
rect 13510 10039 13511 10065
rect 13511 10039 13537 10065
rect 13537 10039 13538 10065
rect 13510 10038 13538 10039
rect 12838 8918 12866 8946
rect 12894 8833 12922 8834
rect 12894 8807 12895 8833
rect 12895 8807 12921 8833
rect 12921 8807 12922 8833
rect 12894 8806 12922 8807
rect 12502 7937 12530 7938
rect 12502 7911 12503 7937
rect 12503 7911 12529 7937
rect 12529 7911 12530 7937
rect 12502 7910 12530 7911
rect 12614 7574 12642 7602
rect 15302 10849 15330 10850
rect 15302 10823 15303 10849
rect 15303 10823 15329 10849
rect 15329 10823 15330 10849
rect 15302 10822 15330 10823
rect 15190 10793 15218 10794
rect 15190 10767 15191 10793
rect 15191 10767 15217 10793
rect 15217 10767 15218 10793
rect 15190 10766 15218 10767
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 13846 10262 13874 10290
rect 14238 10374 14266 10402
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 18830 10598 18858 10626
rect 14910 10401 14938 10402
rect 14910 10375 14911 10401
rect 14911 10375 14937 10401
rect 14937 10375 14938 10401
rect 14910 10374 14938 10375
rect 15022 10345 15050 10346
rect 15022 10319 15023 10345
rect 15023 10319 15049 10345
rect 15049 10319 15050 10345
rect 15022 10318 15050 10319
rect 20006 11102 20034 11130
rect 20006 10766 20034 10794
rect 20006 10457 20034 10458
rect 20006 10431 20007 10457
rect 20007 10431 20033 10457
rect 20033 10431 20034 10457
rect 20006 10430 20034 10431
rect 18942 10318 18970 10346
rect 14350 10289 14378 10290
rect 14350 10263 14351 10289
rect 14351 10263 14377 10289
rect 14377 10263 14378 10289
rect 14350 10262 14378 10263
rect 13846 9617 13874 9618
rect 13846 9591 13847 9617
rect 13847 9591 13873 9617
rect 13873 9591 13874 9617
rect 13846 9590 13874 9591
rect 13734 9534 13762 9562
rect 20006 10038 20034 10066
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 18830 9702 18858 9730
rect 14686 9590 14714 9618
rect 14238 9561 14266 9562
rect 14238 9535 14239 9561
rect 14239 9535 14265 9561
rect 14265 9535 14266 9561
rect 14238 9534 14266 9535
rect 13958 9198 13986 9226
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 20006 9422 20034 9450
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 13398 8918 13426 8946
rect 13286 8806 13314 8834
rect 13566 8862 13594 8890
rect 13398 8750 13426 8778
rect 14294 8889 14322 8890
rect 14294 8863 14295 8889
rect 14295 8863 14321 8889
rect 14321 8863 14322 8889
rect 14294 8862 14322 8863
rect 14630 8833 14658 8834
rect 14630 8807 14631 8833
rect 14631 8807 14657 8833
rect 14657 8807 14658 8833
rect 14630 8806 14658 8807
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 13006 8358 13034 8386
rect 13454 8385 13482 8386
rect 13454 8359 13455 8385
rect 13455 8359 13481 8385
rect 13481 8359 13482 8385
rect 13454 8358 13482 8359
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 12894 7574 12922 7602
rect 13006 7910 13034 7938
rect 13286 7574 13314 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9422 2030 9450 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 10038 2057 10066 2058
rect 10038 2031 10039 2057
rect 10039 2031 10065 2057
rect 10065 2031 10066 2057
rect 10038 2030 10066 2031
rect 10430 1806 10458 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11046 1833 11074 1834
rect 11046 1807 11047 1833
rect 11047 1807 11073 1833
rect 11073 1807 11074 1833
rect 11046 1806 11074 1807
rect 11438 1806 11466 1834
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12446 2030 12474 2058
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9753 18718 9758 18746
rect 9786 18718 10374 18746
rect 10402 18718 10407 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 8745 14238 8750 14266
rect 8778 14238 9366 14266
rect 9394 14238 9399 14266
rect 9473 14238 9478 14266
rect 9506 14238 10150 14266
rect 10178 14238 10183 14266
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 9809 13902 9814 13930
rect 9842 13902 10654 13930
rect 10682 13902 10687 13930
rect 11713 13846 11718 13874
rect 11746 13846 12110 13874
rect 12138 13846 12143 13874
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 10257 13678 10262 13706
rect 10290 13678 11438 13706
rect 11466 13678 11471 13706
rect 9417 13622 9422 13650
rect 9450 13622 10374 13650
rect 10402 13622 11270 13650
rect 11298 13622 11303 13650
rect 8689 13566 8694 13594
rect 8722 13566 9758 13594
rect 9786 13566 9791 13594
rect 11153 13566 11158 13594
rect 11186 13566 11662 13594
rect 11690 13566 11695 13594
rect 2137 13454 2142 13482
rect 2170 13454 5782 13482
rect 5810 13454 7462 13482
rect 7490 13454 7495 13482
rect 10649 13454 10654 13482
rect 10682 13454 10878 13482
rect 10906 13454 12054 13482
rect 12082 13454 12390 13482
rect 12418 13454 12423 13482
rect 11550 13426 11578 13454
rect 7625 13398 7630 13426
rect 7658 13398 10150 13426
rect 10178 13398 11102 13426
rect 11130 13398 11135 13426
rect 11545 13398 11550 13426
rect 11578 13398 11583 13426
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 8129 13230 8134 13258
rect 8162 13230 8862 13258
rect 8890 13230 8895 13258
rect 13449 13174 13454 13202
rect 13482 13174 15974 13202
rect 0 13146 400 13160
rect 15946 13146 15974 13174
rect 20600 13146 21000 13160
rect 0 13118 966 13146
rect 994 13118 999 13146
rect 2137 13118 2142 13146
rect 2170 13118 5726 13146
rect 5754 13118 5759 13146
rect 6841 13118 6846 13146
rect 6874 13118 7798 13146
rect 7826 13118 7831 13146
rect 9641 13118 9646 13146
rect 9674 13118 9679 13146
rect 12889 13118 12894 13146
rect 12922 13118 13342 13146
rect 13370 13118 13375 13146
rect 15946 13118 18830 13146
rect 18858 13118 18863 13146
rect 20113 13118 20118 13146
rect 20146 13118 21000 13146
rect 0 13104 400 13118
rect 7737 13062 7742 13090
rect 7770 13062 8806 13090
rect 8834 13062 8839 13090
rect 9646 13034 9674 13118
rect 20600 13104 21000 13118
rect 7457 13006 7462 13034
rect 7490 13006 9674 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 0 12810 400 12824
rect 20600 12810 21000 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 7401 12782 7406 12810
rect 7434 12782 8190 12810
rect 8218 12782 8223 12810
rect 11489 12782 11494 12810
rect 11522 12782 12782 12810
rect 12810 12782 12815 12810
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 0 12768 400 12782
rect 20600 12768 21000 12782
rect 6897 12726 6902 12754
rect 6930 12726 7350 12754
rect 7378 12726 7383 12754
rect 13449 12726 13454 12754
rect 13482 12726 18830 12754
rect 18858 12726 18863 12754
rect 5721 12670 5726 12698
rect 5754 12670 7854 12698
rect 7882 12670 7887 12698
rect 11601 12670 11606 12698
rect 11634 12670 12390 12698
rect 12418 12670 12423 12698
rect 7345 12614 7350 12642
rect 7378 12614 7910 12642
rect 7938 12614 7943 12642
rect 9249 12614 9254 12642
rect 9282 12614 11550 12642
rect 11578 12614 11583 12642
rect 13426 12614 13678 12642
rect 13706 12614 13711 12642
rect 13393 12558 13398 12586
rect 13426 12558 13454 12614
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 20600 12474 21000 12488
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 20600 12432 21000 12446
rect 9585 12390 9590 12418
rect 9618 12390 11998 12418
rect 12026 12390 12614 12418
rect 12642 12390 12647 12418
rect 12777 12390 12782 12418
rect 12810 12390 18858 12418
rect 18830 12362 18858 12390
rect 8129 12334 8134 12362
rect 8162 12334 10206 12362
rect 10234 12334 10239 12362
rect 11881 12334 11886 12362
rect 11914 12334 12334 12362
rect 12362 12334 12670 12362
rect 12698 12334 15974 12362
rect 18825 12334 18830 12362
rect 18858 12334 18863 12362
rect 15946 12306 15974 12334
rect 15946 12278 18858 12306
rect 18830 12194 18858 12278
rect 18825 12166 18830 12194
rect 18858 12166 18863 12194
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 11265 12110 11270 12138
rect 11298 12110 11550 12138
rect 11578 12110 11583 12138
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 2137 11942 2142 11970
rect 2170 11942 6510 11970
rect 6538 11942 6543 11970
rect 7905 11942 7910 11970
rect 7938 11942 10654 11970
rect 10682 11942 11158 11970
rect 11186 11942 11191 11970
rect 8073 11830 8078 11858
rect 8106 11830 8470 11858
rect 8498 11830 8503 11858
rect 11489 11830 11494 11858
rect 11522 11830 11942 11858
rect 11970 11830 11975 11858
rect 0 11802 400 11816
rect 20600 11802 21000 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 10817 11774 10822 11802
rect 10850 11774 11270 11802
rect 11298 11774 11303 11802
rect 12441 11774 12446 11802
rect 12474 11774 13146 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 7009 11718 7014 11746
rect 7042 11718 7462 11746
rect 7490 11718 7495 11746
rect 8185 11718 8190 11746
rect 8218 11718 8694 11746
rect 8722 11718 8727 11746
rect 10369 11718 10374 11746
rect 10402 11718 10766 11746
rect 10794 11718 10799 11746
rect 13118 11690 13146 11774
rect 20600 11760 21000 11774
rect 13113 11662 13118 11690
rect 13146 11662 13398 11690
rect 13426 11662 14798 11690
rect 14826 11662 14831 11690
rect 7569 11606 7574 11634
rect 7602 11606 8190 11634
rect 8218 11606 8223 11634
rect 10033 11606 10038 11634
rect 10066 11606 10318 11634
rect 10346 11606 10351 11634
rect 2137 11550 2142 11578
rect 2170 11550 4214 11578
rect 8409 11550 8414 11578
rect 8442 11550 8862 11578
rect 8890 11550 9254 11578
rect 9282 11550 9287 11578
rect 10089 11550 10094 11578
rect 10122 11550 10654 11578
rect 10682 11550 10687 11578
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 4186 11522 4214 11550
rect 15946 11522 15974 11550
rect 4186 11494 4942 11522
rect 4970 11494 6286 11522
rect 6314 11494 6319 11522
rect 7513 11494 7518 11522
rect 7546 11494 9590 11522
rect 9618 11494 10794 11522
rect 13785 11494 13790 11522
rect 13818 11494 14574 11522
rect 14602 11494 15974 11522
rect 0 11466 400 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 0 11424 400 11438
rect 10766 11410 10794 11494
rect 20600 11466 21000 11480
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 10761 11382 10766 11410
rect 10794 11382 11550 11410
rect 11578 11382 11583 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 8689 11214 8694 11242
rect 8722 11214 13174 11242
rect 13202 11214 13207 11242
rect 7793 11158 7798 11186
rect 7826 11158 8078 11186
rect 8106 11158 8750 11186
rect 8778 11158 8783 11186
rect 9305 11158 9310 11186
rect 9338 11158 10094 11186
rect 10122 11158 10127 11186
rect 10859 11158 10878 11186
rect 10906 11158 10911 11186
rect 20600 11130 21000 11144
rect 6505 11102 6510 11130
rect 6538 11102 8190 11130
rect 8218 11102 8223 11130
rect 9025 11102 9030 11130
rect 9058 11102 9422 11130
rect 9450 11102 11606 11130
rect 11634 11102 11639 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 2081 11046 2086 11074
rect 2114 11046 9086 11074
rect 9114 11046 9534 11074
rect 9562 11046 9567 11074
rect 13169 11046 13174 11074
rect 13202 11046 13678 11074
rect 13706 11046 13711 11074
rect 7009 10990 7014 11018
rect 7042 10990 9590 11018
rect 9618 10990 9623 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 6286 10934 6342 10962
rect 6370 10934 6790 10962
rect 6818 10934 7406 10962
rect 7434 10934 7910 10962
rect 7938 10934 7943 10962
rect 8073 10934 8078 10962
rect 8106 10934 8246 10962
rect 8274 10934 8279 10962
rect 10369 10934 10374 10962
rect 10402 10934 10766 10962
rect 10794 10934 11158 10962
rect 11186 10934 11191 10962
rect 6286 10906 6314 10934
rect 5329 10878 5334 10906
rect 5362 10878 6314 10906
rect 6734 10878 7350 10906
rect 7378 10878 7383 10906
rect 10929 10878 10934 10906
rect 10962 10878 11438 10906
rect 11466 10878 11471 10906
rect 13113 10878 13118 10906
rect 13146 10878 13342 10906
rect 13370 10878 13566 10906
rect 13594 10878 13599 10906
rect 6734 10850 6762 10878
rect 6001 10822 6006 10850
rect 6034 10822 6762 10850
rect 7177 10822 7182 10850
rect 7210 10822 11326 10850
rect 11354 10822 11359 10850
rect 15297 10822 15302 10850
rect 15330 10822 18858 10850
rect 18830 10794 18858 10822
rect 20600 10794 21000 10808
rect 6393 10766 6398 10794
rect 6426 10766 6958 10794
rect 6986 10766 6991 10794
rect 7289 10766 7294 10794
rect 7322 10766 7574 10794
rect 7602 10766 7607 10794
rect 8017 10766 8022 10794
rect 8050 10766 8302 10794
rect 8330 10766 8694 10794
rect 8722 10766 8727 10794
rect 9193 10766 9198 10794
rect 9226 10766 11662 10794
rect 11690 10766 11695 10794
rect 15185 10766 15190 10794
rect 15218 10766 15974 10794
rect 18825 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 5665 10710 5670 10738
rect 5698 10710 7686 10738
rect 7714 10710 7719 10738
rect 7905 10710 7910 10738
rect 7938 10710 9254 10738
rect 9282 10710 13398 10738
rect 13426 10710 13431 10738
rect 15946 10682 15974 10766
rect 20600 10752 21000 10766
rect 6729 10654 6734 10682
rect 6762 10654 8470 10682
rect 8498 10654 8862 10682
rect 8890 10654 8895 10682
rect 15946 10654 18858 10682
rect 18830 10626 18858 10654
rect 18825 10598 18830 10626
rect 18858 10598 18863 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 10201 10542 10206 10570
rect 10234 10542 10934 10570
rect 10962 10542 10967 10570
rect 20600 10458 21000 10472
rect 6841 10430 6846 10458
rect 6874 10430 7742 10458
rect 7770 10430 7775 10458
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 20600 10416 21000 10430
rect 10033 10374 10038 10402
rect 10066 10374 11382 10402
rect 11410 10374 11415 10402
rect 14233 10374 14238 10402
rect 14266 10374 14910 10402
rect 14938 10374 14943 10402
rect 9137 10318 9142 10346
rect 9170 10318 10766 10346
rect 10794 10318 10799 10346
rect 15017 10318 15022 10346
rect 15050 10318 18942 10346
rect 18970 10318 18975 10346
rect 9254 10262 10654 10290
rect 10682 10262 10687 10290
rect 13841 10262 13846 10290
rect 13874 10262 14350 10290
rect 14378 10262 14383 10290
rect 9254 10234 9282 10262
rect 7401 10206 7406 10234
rect 7434 10206 8078 10234
rect 8106 10206 8526 10234
rect 8554 10206 8559 10234
rect 9249 10206 9254 10234
rect 9282 10206 9287 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 7457 10150 7462 10178
rect 7490 10150 7495 10178
rect 7462 10066 7490 10150
rect 20600 10122 21000 10136
rect 8185 10094 8190 10122
rect 8218 10094 9618 10122
rect 10033 10094 10038 10122
rect 10066 10094 11102 10122
rect 11130 10094 13622 10122
rect 13650 10094 13655 10122
rect 20006 10094 21000 10122
rect 9590 10066 9618 10094
rect 20006 10066 20034 10094
rect 20600 10080 21000 10094
rect 7462 10038 7966 10066
rect 7994 10038 8414 10066
rect 8442 10038 8447 10066
rect 9585 10038 9590 10066
rect 9618 10038 9623 10066
rect 9809 10038 9814 10066
rect 9842 10038 10878 10066
rect 10906 10038 10911 10066
rect 12721 10038 12726 10066
rect 12754 10038 13230 10066
rect 13258 10038 13263 10066
rect 13426 10038 13510 10066
rect 13538 10038 13543 10066
rect 20001 10038 20006 10066
rect 20034 10038 20039 10066
rect 13426 10010 13454 10038
rect 4993 9982 4998 10010
rect 5026 9982 7126 10010
rect 7154 9982 7159 10010
rect 8353 9982 8358 10010
rect 8386 9982 9366 10010
rect 9394 9982 9399 10010
rect 9977 9982 9982 10010
rect 10010 9982 10262 10010
rect 10290 9982 10295 10010
rect 11209 9982 11214 10010
rect 11242 9982 12838 10010
rect 12866 9982 13454 10010
rect 8969 9926 8974 9954
rect 9002 9926 9534 9954
rect 9562 9926 9567 9954
rect 11041 9926 11046 9954
rect 11074 9926 11494 9954
rect 11522 9926 11662 9954
rect 11690 9926 11695 9954
rect 12161 9926 12166 9954
rect 12194 9926 12670 9954
rect 12698 9926 12703 9954
rect 7401 9870 7406 9898
rect 7434 9870 7490 9898
rect 10985 9870 10990 9898
rect 11018 9870 11550 9898
rect 11578 9870 11583 9898
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 7462 9674 7490 9870
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 8857 9702 8862 9730
rect 8890 9702 12782 9730
rect 12810 9702 12815 9730
rect 15946 9702 18830 9730
rect 18858 9702 18863 9730
rect 15946 9674 15974 9702
rect 4186 9646 4998 9674
rect 5026 9646 5031 9674
rect 7457 9646 7462 9674
rect 7490 9646 7495 9674
rect 10990 9646 11326 9674
rect 11354 9646 11718 9674
rect 11746 9646 11751 9674
rect 13225 9646 13230 9674
rect 13258 9646 15974 9674
rect 4186 9618 4214 9646
rect 10990 9618 11018 9646
rect 2137 9590 2142 9618
rect 2170 9590 4214 9618
rect 6449 9590 6454 9618
rect 6482 9590 6790 9618
rect 6818 9590 6823 9618
rect 7233 9590 7238 9618
rect 7266 9590 7630 9618
rect 7658 9590 7663 9618
rect 7961 9590 7966 9618
rect 7994 9590 9086 9618
rect 9114 9590 9119 9618
rect 9193 9590 9198 9618
rect 9226 9590 10654 9618
rect 10682 9590 10687 9618
rect 10985 9590 10990 9618
rect 11018 9590 11023 9618
rect 13841 9590 13846 9618
rect 13874 9590 14686 9618
rect 14714 9590 18830 9618
rect 18858 9590 18863 9618
rect 6729 9534 6734 9562
rect 6762 9534 7126 9562
rect 7154 9534 7742 9562
rect 7770 9534 7775 9562
rect 8297 9534 8302 9562
rect 8330 9534 9422 9562
rect 9450 9534 10822 9562
rect 10850 9534 12558 9562
rect 12586 9534 12591 9562
rect 13729 9534 13734 9562
rect 13762 9534 14238 9562
rect 14266 9534 14271 9562
rect 7345 9478 7350 9506
rect 7378 9478 9758 9506
rect 9786 9478 10038 9506
rect 10066 9478 10071 9506
rect 0 9450 400 9464
rect 20600 9450 21000 9464
rect 0 9422 966 9450
rect 994 9422 999 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 0 9408 400 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 6057 9310 6062 9338
rect 6090 9310 7126 9338
rect 7154 9310 7159 9338
rect 10761 9310 10766 9338
rect 10794 9310 10878 9338
rect 10906 9310 10911 9338
rect 7513 9254 7518 9282
rect 7546 9254 8918 9282
rect 8946 9254 8951 9282
rect 6953 9198 6958 9226
rect 6986 9198 7462 9226
rect 7490 9198 7495 9226
rect 8129 9198 8134 9226
rect 8162 9198 8414 9226
rect 8442 9198 8447 9226
rect 8969 9198 8974 9226
rect 9002 9198 9814 9226
rect 9842 9198 9847 9226
rect 10593 9198 10598 9226
rect 10626 9198 11270 9226
rect 11298 9198 11303 9226
rect 11657 9198 11662 9226
rect 11690 9198 11886 9226
rect 11914 9198 13958 9226
rect 13986 9198 13991 9226
rect 6897 9142 6902 9170
rect 6930 9142 8246 9170
rect 8274 9142 8279 9170
rect 8974 9114 9002 9198
rect 10089 9142 10094 9170
rect 10122 9142 10822 9170
rect 10850 9142 11718 9170
rect 11746 9142 11751 9170
rect 11825 9142 11830 9170
rect 11858 9142 12334 9170
rect 12362 9142 12367 9170
rect 6673 9086 6678 9114
rect 6706 9086 7238 9114
rect 7266 9086 8078 9114
rect 8106 9086 8111 9114
rect 8185 9086 8190 9114
rect 8218 9086 9002 9114
rect 7177 9030 7182 9058
rect 7210 9030 10206 9058
rect 10234 9030 10239 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 7961 8918 7966 8946
rect 7994 8918 10598 8946
rect 10626 8918 10631 8946
rect 11881 8918 11886 8946
rect 11914 8918 12838 8946
rect 12866 8918 13398 8946
rect 13426 8918 13431 8946
rect 13561 8862 13566 8890
rect 13594 8862 14294 8890
rect 14322 8862 15974 8890
rect 15946 8834 15974 8862
rect 8241 8806 8246 8834
rect 8274 8806 8582 8834
rect 8610 8806 8615 8834
rect 9697 8806 9702 8834
rect 9730 8806 11858 8834
rect 12329 8806 12334 8834
rect 12362 8806 12894 8834
rect 12922 8806 13286 8834
rect 13314 8806 14630 8834
rect 14658 8806 14663 8834
rect 15946 8806 18830 8834
rect 18858 8806 18863 8834
rect 11830 8778 11858 8806
rect 20600 8778 21000 8792
rect 11214 8750 11718 8778
rect 11746 8750 11751 8778
rect 11830 8750 11998 8778
rect 12026 8750 13398 8778
rect 13426 8750 13431 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 11214 8722 11242 8750
rect 20600 8736 21000 8750
rect 7849 8694 7854 8722
rect 7882 8694 11214 8722
rect 11242 8694 11247 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 10761 8582 10766 8610
rect 10794 8582 11550 8610
rect 11578 8582 11583 8610
rect 8801 8526 8806 8554
rect 8834 8526 9310 8554
rect 9338 8526 9926 8554
rect 9954 8526 9959 8554
rect 11153 8526 11158 8554
rect 11186 8526 11606 8554
rect 11634 8526 11639 8554
rect 5833 8470 5838 8498
rect 5866 8470 6958 8498
rect 6986 8470 9254 8498
rect 9282 8470 9814 8498
rect 9842 8470 9982 8498
rect 10010 8470 10015 8498
rect 10593 8470 10598 8498
rect 10626 8470 11662 8498
rect 11690 8470 11695 8498
rect 5497 8414 5502 8442
rect 5530 8414 5535 8442
rect 6897 8414 6902 8442
rect 6930 8414 7350 8442
rect 7378 8414 7574 8442
rect 7602 8414 7607 8442
rect 7686 8414 7798 8442
rect 7826 8414 7831 8442
rect 9025 8414 9030 8442
rect 9058 8414 10430 8442
rect 10458 8414 10463 8442
rect 11209 8414 11214 8442
rect 11242 8414 11802 8442
rect 5502 8386 5530 8414
rect 7686 8386 7714 8414
rect 5502 8358 6342 8386
rect 6370 8358 6790 8386
rect 6818 8358 6823 8386
rect 7625 8358 7630 8386
rect 7658 8358 7714 8386
rect 10033 8358 10038 8386
rect 10066 8358 10934 8386
rect 10962 8358 10967 8386
rect 11774 8330 11802 8414
rect 13001 8358 13006 8386
rect 13034 8358 13454 8386
rect 13482 8358 13487 8386
rect 9585 8302 9590 8330
rect 9618 8302 10598 8330
rect 10626 8302 10631 8330
rect 11769 8302 11774 8330
rect 11802 8302 11807 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 7737 8134 7742 8162
rect 7770 8134 8694 8162
rect 8722 8134 8727 8162
rect 9361 8134 9366 8162
rect 9394 8134 9534 8162
rect 9562 8134 9567 8162
rect 9809 8134 9814 8162
rect 9842 8134 11046 8162
rect 11074 8134 11326 8162
rect 11354 8134 11359 8162
rect 8801 7966 8806 7994
rect 8834 7966 9590 7994
rect 9618 7966 9623 7994
rect 11321 7966 11326 7994
rect 11354 7966 12110 7994
rect 12138 7966 12143 7994
rect 6673 7910 6678 7938
rect 6706 7910 7686 7938
rect 7714 7910 7719 7938
rect 9305 7910 9310 7938
rect 9338 7910 10206 7938
rect 10234 7910 10239 7938
rect 12497 7910 12502 7938
rect 12530 7910 13006 7938
rect 13034 7910 13039 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 7681 7686 7686 7714
rect 7714 7686 9142 7714
rect 9170 7686 9175 7714
rect 9473 7686 9478 7714
rect 9506 7686 10374 7714
rect 10402 7686 10407 7714
rect 9529 7630 9534 7658
rect 9562 7630 10206 7658
rect 10234 7630 11606 7658
rect 11634 7630 11639 7658
rect 6337 7574 6342 7602
rect 6370 7574 7014 7602
rect 7042 7574 7350 7602
rect 7378 7574 7966 7602
rect 7994 7574 8750 7602
rect 8778 7574 8783 7602
rect 11545 7574 11550 7602
rect 11578 7574 12614 7602
rect 12642 7574 12894 7602
rect 12922 7574 13286 7602
rect 13314 7574 13319 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 8857 7350 8862 7378
rect 8890 7350 8895 7378
rect 8862 7322 8890 7350
rect 8745 7294 8750 7322
rect 8778 7294 9534 7322
rect 9562 7294 9567 7322
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 9417 2030 9422 2058
rect 9450 2030 10038 2058
rect 10066 2030 10071 2058
rect 12441 2030 12446 2058
rect 12474 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10425 1806 10430 1834
rect 10458 1806 11046 1834
rect 11074 1806 11079 1834
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 10878 11158 10906 11186
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 10878 9310 10906 9338
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 10878 11186 10906 11191
rect 10878 9338 10906 11158
rect 10878 9305 10906 9310
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7504 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6608 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7224 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _103_
timestamp 1698175906
transform 1 0 8008 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1698175906
transform 1 0 8512 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform 1 0 8792 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11648 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _107_
timestamp 1698175906
transform -1 0 10080 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _108_
timestamp 1698175906
transform -1 0 9968 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10864 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform 1 0 10080 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform -1 0 10920 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7560 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform 1 0 10528 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 11536 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10808 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _116_
timestamp 1698175906
transform 1 0 6832 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 7672 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _118_
timestamp 1698175906
transform -1 0 8568 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 9016 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 9968 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10584 0 -1 7840
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _122_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 7840
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8064 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9464 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 7840 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 11648 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _127_
timestamp 1698175906
transform 1 0 13608 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _128_
timestamp 1698175906
transform -1 0 13608 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform -1 0 7560 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 9520 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform 1 0 10584 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform -1 0 9352 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform -1 0 9520 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9072 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8344 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform -1 0 8512 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _139_
timestamp 1698175906
transform -1 0 7840 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform 1 0 8288 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform 1 0 10136 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _142_
timestamp 1698175906
transform -1 0 9464 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9016 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _144_
timestamp 1698175906
transform 1 0 8680 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 6944 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _146_
timestamp 1698175906
transform 1 0 7560 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 8344 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _149_
timestamp 1698175906
transform -1 0 8400 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _150_
timestamp 1698175906
transform 1 0 8064 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _151_
timestamp 1698175906
transform 1 0 11648 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _152_
timestamp 1698175906
transform 1 0 13664 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _153_
timestamp 1698175906
transform -1 0 13664 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 1 10192
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _156_
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform -1 0 10920 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 8008 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7728 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform -1 0 9856 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _161_
timestamp 1698175906
transform 1 0 13328 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13160 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7616 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _164_
timestamp 1698175906
transform -1 0 7672 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _165_
timestamp 1698175906
transform -1 0 7560 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _166_
timestamp 1698175906
transform -1 0 7616 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform -1 0 10192 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11480 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 -1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _170_
timestamp 1698175906
transform -1 0 10192 0 -1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform 1 0 14112 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _172_
timestamp 1698175906
transform -1 0 13888 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 12656 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _174_
timestamp 1698175906
transform -1 0 11928 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _175_
timestamp 1698175906
transform -1 0 12376 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _176_
timestamp 1698175906
transform -1 0 9632 0 -1 8624
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _177_
timestamp 1698175906
transform 1 0 8624 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9744 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _179_
timestamp 1698175906
transform 1 0 9016 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10360 0 1 10976
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _181_
timestamp 1698175906
transform -1 0 9800 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _182_
timestamp 1698175906
transform 1 0 9296 0 1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform -1 0 9632 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform 1 0 9912 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _185_
timestamp 1698175906
transform -1 0 11536 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _186_
timestamp 1698175906
transform -1 0 12096 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _187_
timestamp 1698175906
transform 1 0 10976 0 1 11760
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _188_
timestamp 1698175906
transform -1 0 7560 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11984 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _190_
timestamp 1698175906
transform 1 0 7336 0 -1 13328
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_
timestamp 1698175906
transform 1 0 6216 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _192_
timestamp 1698175906
transform 1 0 6888 0 -1 10976
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1698175906
transform 1 0 12656 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _194_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _195_
timestamp 1698175906
transform -1 0 11592 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11088 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _197_
timestamp 1698175906
transform -1 0 10472 0 1 13328
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _198_
timestamp 1698175906
transform -1 0 11816 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _199_
timestamp 1698175906
transform -1 0 11368 0 1 13328
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8848 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 13048 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform 1 0 7672 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 5376 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 6216 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 8400 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 5208 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform -1 0 8064 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 13160 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 11704 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform -1 0 7280 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 12768 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform -1 0 6552 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 10808 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 13440 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 11480 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 7224 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 10808 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform -1 0 7336 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform -1 0 6496 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 11928 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 9800 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 10584 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _226_
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _227_
timestamp 1698175906
transform 1 0 14784 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _228_
timestamp 1698175906
transform 1 0 13216 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _229_
timestamp 1698175906
transform 1 0 15064 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13160 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__A3
timestamp 1698175906
transform 1 0 8680 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__A2
timestamp 1698175906
transform 1 0 14224 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__A1
timestamp 1698175906
transform -1 0 8232 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 9744 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 7000 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 7952 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 10192 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 6832 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 8064 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 13328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 7392 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 14616 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 6776 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 13328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform -1 0 13328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform -1 0 8960 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform -1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 12432 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 8120 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 6776 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 13664 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 11536 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform -1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9072 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9464 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10360 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11312 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_154 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9296 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_162 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 11928 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 12040 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 9072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 9408 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183
timestamp 1698175906
transform 1 0 10920 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 11816 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_148
timestamp 1698175906
transform 1 0 8960 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_180
timestamp 1698175906
transform 1 0 10752 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_196
timestamp 1698175906
transform 1 0 11648 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_204
timestamp 1698175906
transform 1 0 12096 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_222
timestamp 1698175906
transform 1 0 13104 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_226
timestamp 1698175906
transform 1 0 13328 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 14224 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_88
timestamp 1698175906
transform 1 0 5600 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_96
timestamp 1698175906
transform 1 0 6048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_98
timestamp 1698175906
transform 1 0 6160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_128
timestamp 1698175906
transform 1 0 7840 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_132
timestamp 1698175906
transform 1 0 8064 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 8848 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_148
timestamp 1698175906
transform 1 0 8960 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_157
timestamp 1698175906
transform 1 0 9464 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_165
timestamp 1698175906
transform 1 0 9912 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_177
timestamp 1698175906
transform 1 0 10584 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_216
timestamp 1698175906
transform 1 0 12768 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698175906
transform 1 0 6888 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698175906
transform 1 0 7112 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698175906
transform 1 0 7336 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_121
timestamp 1698175906
transform 1 0 7448 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_128
timestamp 1698175906
transform 1 0 7840 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_136
timestamp 1698175906
transform 1 0 8288 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_140
timestamp 1698175906
transform 1 0 8512 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_214
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_230
timestamp 1698175906
transform 1 0 13552 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_238
timestamp 1698175906
transform 1 0 14000 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 5152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_113
timestamp 1698175906
transform 1 0 7000 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_115
timestamp 1698175906
transform 1 0 7112 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_122
timestamp 1698175906
transform 1 0 7504 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 8344 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698175906
transform 1 0 9072 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_152
timestamp 1698175906
transform 1 0 9184 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_160
timestamp 1698175906
transform 1 0 9632 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_170
timestamp 1698175906
transform 1 0 10192 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_172
timestamp 1698175906
transform 1 0 10304 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_203
timestamp 1698175906
transform 1 0 12040 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698175906
transform 1 0 12992 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_224
timestamp 1698175906
transform 1 0 13216 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_232
timestamp 1698175906
transform 1 0 13664 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_264
timestamp 1698175906
transform 1 0 15456 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_131
timestamp 1698175906
transform 1 0 8008 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_146
timestamp 1698175906
transform 1 0 8848 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_162
timestamp 1698175906
transform 1 0 9744 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698175906
transform 1 0 10192 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_183
timestamp 1698175906
transform 1 0 10920 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_191
timestamp 1698175906
transform 1 0 11368 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_195
timestamp 1698175906
transform 1 0 11592 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_202
timestamp 1698175906
transform 1 0 11984 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_210
timestamp 1698175906
transform 1 0 12432 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_214
timestamp 1698175906
transform 1 0 12656 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 14728 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_104
timestamp 1698175906
transform 1 0 6496 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_124
timestamp 1698175906
transform 1 0 7616 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_126
timestamp 1698175906
transform 1 0 7728 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698175906
transform 1 0 8344 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_150
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_172
timestamp 1698175906
transform 1 0 10304 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_187
timestamp 1698175906
transform 1 0 11144 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_195
timestamp 1698175906
transform 1 0 11592 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_202
timestamp 1698175906
transform 1 0 11984 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698175906
transform 1 0 12656 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_252
timestamp 1698175906
transform 1 0 14784 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_268
timestamp 1698175906
transform 1 0 15680 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 16128 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 4760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 4872 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 6888 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_155
timestamp 1698175906
transform 1 0 9352 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_163
timestamp 1698175906
transform 1 0 9800 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_170
timestamp 1698175906
transform 1 0 10192 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_183
timestamp 1698175906
transform 1 0 10920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_187
timestamp 1698175906
transform 1 0 11144 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_196
timestamp 1698175906
transform 1 0 11648 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_240
timestamp 1698175906
transform 1 0 14112 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_112
timestamp 1698175906
transform 1 0 6944 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_124
timestamp 1698175906
transform 1 0 7616 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_146
timestamp 1698175906
transform 1 0 8848 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_202
timestamp 1698175906
transform 1 0 11984 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_220
timestamp 1698175906
transform 1 0 12992 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_224
timestamp 1698175906
transform 1 0 13216 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_236
timestamp 1698175906
transform 1 0 13888 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_268
timestamp 1698175906
transform 1 0 15680 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 16128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698175906
transform 1 0 6776 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 10360 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_251
timestamp 1698175906
transform 1 0 14728 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_258
timestamp 1698175906
transform 1 0 15120 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_290
timestamp 1698175906
transform 1 0 16912 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_306
timestamp 1698175906
transform 1 0 17808 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698175906
transform 1 0 18256 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_80
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_110
timestamp 1698175906
transform 1 0 6832 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 8400 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 12264 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_217
timestamp 1698175906
transform 1 0 12824 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_225
timestamp 1698175906
transform 1 0 13272 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_263
timestamp 1698175906
transform 1 0 15400 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 4536 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 4760 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698175906
transform 1 0 6496 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_111
timestamp 1698175906
transform 1 0 6888 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_127
timestamp 1698175906
transform 1 0 7784 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_131
timestamp 1698175906
transform 1 0 8008 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_141
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_145
timestamp 1698175906
transform 1 0 8792 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_149
timestamp 1698175906
transform 1 0 9016 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698175906
transform 1 0 10360 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_200
timestamp 1698175906
transform 1 0 11872 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_216
timestamp 1698175906
transform 1 0 12768 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_220
timestamp 1698175906
transform 1 0 12992 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_222
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_239
timestamp 1698175906
transform 1 0 14056 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_96
timestamp 1698175906
transform 1 0 6048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_98
timestamp 1698175906
transform 1 0 6160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_151
timestamp 1698175906
transform 1 0 9128 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_166
timestamp 1698175906
transform 1 0 9968 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_174
timestamp 1698175906
transform 1 0 10416 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_176
timestamp 1698175906
transform 1 0 10528 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_183
timestamp 1698175906
transform 1 0 10920 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_199
timestamp 1698175906
transform 1 0 11816 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 12264 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_220
timestamp 1698175906
transform 1 0 12992 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_250
timestamp 1698175906
transform 1 0 14672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_254
timestamp 1698175906
transform 1 0 14896 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_270
timestamp 1698175906
transform 1 0 15792 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 16240 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698175906
transform 1 0 7560 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_131
timestamp 1698175906
transform 1 0 8008 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_134
timestamp 1698175906
transform 1 0 8176 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698175906
transform 1 0 10024 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_183
timestamp 1698175906
transform 1 0 10920 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_204
timestamp 1698175906
transform 1 0 12096 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_208
timestamp 1698175906
transform 1 0 12320 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_212
timestamp 1698175906
transform 1 0 12544 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_118
timestamp 1698175906
transform 1 0 7280 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_122
timestamp 1698175906
transform 1 0 7504 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_168
timestamp 1698175906
transform 1 0 10080 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_172
timestamp 1698175906
transform 1 0 10304 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_180
timestamp 1698175906
transform 1 0 10752 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_218
timestamp 1698175906
transform 1 0 12880 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_250
timestamp 1698175906
transform 1 0 14672 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698175906
transform 1 0 15568 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 16016 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_115
timestamp 1698175906
transform 1 0 7112 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_131
timestamp 1698175906
transform 1 0 8008 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_135
timestamp 1698175906
transform 1 0 8232 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_167
timestamp 1698175906
transform 1 0 10024 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_199
timestamp 1698175906
transform 1 0 11816 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_230
timestamp 1698175906
transform 1 0 13552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_234
timestamp 1698175906
transform 1 0 13776 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_131
timestamp 1698175906
transform 1 0 8008 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_135
timestamp 1698175906
transform 1 0 8232 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_155
timestamp 1698175906
transform 1 0 9352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_192
timestamp 1698175906
transform 1 0 11424 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_196
timestamp 1698175906
transform 1 0 11648 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_204
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_220
timestamp 1698175906
transform 1 0 12992 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_230
timestamp 1698175906
transform 1 0 13552 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_262
timestamp 1698175906
transform 1 0 15344 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 16240 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 2240 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 2464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_115
timestamp 1698175906
transform 1 0 7112 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_160
timestamp 1698175906
transform 1 0 9632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_164
timestamp 1698175906
transform 1 0 9856 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_199
timestamp 1698175906
transform 1 0 11816 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_231
timestamp 1698175906
transform 1 0 13608 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698175906
transform 1 0 14056 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 14280 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_333
timestamp 1698175906
transform 1 0 19320 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_341
timestamp 1698175906
transform 1 0 19768 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_171
timestamp 1698175906
transform 1 0 10248 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_175
timestamp 1698175906
transform 1 0 10472 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_139
timestamp 1698175906
transform 1 0 8456 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_147
timestamp 1698175906
transform 1 0 8904 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_151
timestamp 1698175906
transform 1 0 9128 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_153
timestamp 1698175906
transform 1 0 9240 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_160
timestamp 1698175906
transform 1 0 9632 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_168
timestamp 1698175906
transform 1 0 10080 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 10304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 10416 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698175906
transform 1 0 9520 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 9744 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_189
timestamp 1698175906
transform 1 0 11256 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698175906
transform 1 0 12152 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita6_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita6_26
timestamp 1698175906
transform 1 0 9968 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2240 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 12096 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 2240 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 9464 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 9800 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 10472 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 9408 400 9464 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 6692 7812 6692 7812 0 _000_
rlabel metal2 8848 11676 8848 11676 0 _001_
rlabel metal3 6692 10724 6692 10724 0 _002_
rlabel metal3 7896 11620 7896 11620 0 _003_
rlabel metal2 13636 9296 13636 9296 0 _004_
rlabel metal2 12180 9800 12180 9800 0 _005_
rlabel metal2 6804 12572 6804 12572 0 _006_
rlabel metal2 13244 9100 13244 9100 0 _007_
rlabel metal2 6076 9436 6076 9436 0 _008_
rlabel metal2 11284 8064 11284 8064 0 _009_
rlabel metal2 13748 10416 13748 10416 0 _010_
rlabel metal2 11956 7420 11956 7420 0 _011_
rlabel metal3 8428 7700 8428 7700 0 _012_
rlabel metal2 9380 13748 9380 13748 0 _013_
rlabel metal2 11396 12152 11396 12152 0 _014_
rlabel metal3 7336 13132 7336 13132 0 _015_
rlabel metal3 7056 10892 7056 10892 0 _016_
rlabel metal3 12012 12684 12012 12684 0 _017_
rlabel metal2 10332 13300 10332 13300 0 _018_
rlabel metal2 11088 13580 11088 13580 0 _019_
rlabel metal3 9772 7924 9772 7924 0 _020_
rlabel metal2 13468 11368 13468 11368 0 _021_
rlabel metal3 8512 13244 8512 13244 0 _022_
rlabel metal2 6972 8596 6972 8596 0 _023_
rlabel metal2 12852 9016 12852 9016 0 _024_
rlabel metal2 13804 9464 13804 9464 0 _025_
rlabel metal2 12656 10052 12656 10052 0 _026_
rlabel metal3 13482 10052 13482 10052 0 _027_
rlabel metal2 10668 11928 10668 11928 0 _028_
rlabel metal2 7700 12684 7700 12684 0 _029_
rlabel metal2 9632 8428 9632 8428 0 _030_
rlabel metal2 13020 8736 13020 8736 0 _031_
rlabel metal2 7336 9716 7336 9716 0 _032_
rlabel metal2 7364 9212 7364 9212 0 _033_
rlabel metal2 7252 9352 7252 9352 0 _034_
rlabel metal3 10500 8372 10500 8372 0 _035_
rlabel metal2 11116 8512 11116 8512 0 _036_
rlabel metal2 10976 13468 10976 13468 0 _037_
rlabel metal3 14112 10276 14112 10276 0 _038_
rlabel metal2 12348 7980 12348 7980 0 _039_
rlabel metal2 12012 7952 12012 7952 0 _040_
rlabel metal2 9268 8008 9268 8008 0 _041_
rlabel metal2 9100 7896 9100 7896 0 _042_
rlabel metal2 9380 7812 9380 7812 0 _043_
rlabel metal2 7476 12376 7476 12376 0 _044_
rlabel metal2 10388 13580 10388 13580 0 _045_
rlabel metal2 9548 14000 9548 14000 0 _046_
rlabel metal2 10948 10864 10948 10864 0 _047_
rlabel metal2 11424 11900 11424 11900 0 _048_
rlabel metal3 11732 11844 11732 11844 0 _049_
rlabel metal2 7420 13272 7420 13272 0 _050_
rlabel metal2 11172 12180 11172 12180 0 _051_
rlabel metal3 6692 10780 6692 10780 0 _052_
rlabel metal2 11508 12768 11508 12768 0 _053_
rlabel metal2 10276 13580 10276 13580 0 _054_
rlabel metal2 10332 12460 10332 12460 0 _055_
rlabel metal2 11172 13524 11172 13524 0 _056_
rlabel metal2 7252 8820 7252 8820 0 _057_
rlabel metal2 6748 9380 6748 9380 0 _058_
rlabel metal2 8260 9044 8260 9044 0 _059_
rlabel metal2 8792 8764 8792 8764 0 _060_
rlabel metal2 11032 10388 11032 10388 0 _061_
rlabel metal2 11900 8624 11900 8624 0 _062_
rlabel metal2 9828 11592 9828 11592 0 _063_
rlabel metal2 7532 10780 7532 10780 0 _064_
rlabel metal2 11340 8288 11340 8288 0 _065_
rlabel metal2 10836 8988 10836 8988 0 _066_
rlabel metal2 9604 8008 9604 8008 0 _067_
rlabel metal2 10612 9072 10612 9072 0 _068_
rlabel metal2 10976 11956 10976 11956 0 _069_
rlabel metal3 9744 8428 9744 8428 0 _070_
rlabel metal2 10164 8092 10164 8092 0 _071_
rlabel metal2 7476 9184 7476 9184 0 _072_
rlabel metal3 9604 10080 9604 10080 0 _073_
rlabel metal2 7476 10220 7476 10220 0 _074_
rlabel metal2 9268 9884 9268 9884 0 _075_
rlabel metal2 7028 10206 7028 10206 0 _076_
rlabel metal2 10332 7812 10332 7812 0 _077_
rlabel metal2 8372 9548 8372 9548 0 _078_
rlabel metal3 11340 10724 11340 10724 0 _079_
rlabel metal2 13776 9604 13776 9604 0 _080_
rlabel metal2 14196 10780 14196 10780 0 _081_
rlabel metal2 13636 11172 13636 11172 0 _082_
rlabel metal2 9996 9800 9996 9800 0 _083_
rlabel metal2 7084 10220 7084 10220 0 _084_
rlabel metal2 7588 12600 7588 12600 0 _085_
rlabel metal2 9212 9800 9212 9800 0 _086_
rlabel metal2 11284 11872 11284 11872 0 _087_
rlabel metal2 9100 13160 9100 13160 0 _088_
rlabel metal3 9072 14252 9072 14252 0 _089_
rlabel metal2 7644 8176 7644 8176 0 _090_
rlabel metal2 7812 11004 7812 11004 0 _091_
rlabel metal2 7420 10500 7420 10500 0 _092_
rlabel metal2 10780 10360 10780 10360 0 _093_
rlabel metal2 8932 9408 8932 9408 0 _094_
rlabel metal3 10836 9716 10836 9716 0 _095_
rlabel metal2 7308 10584 7308 10584 0 _096_
rlabel metal2 9436 9044 9436 9044 0 _097_
rlabel metal2 8232 11284 8232 11284 0 _098_
rlabel metal2 8148 11144 8148 11144 0 _099_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal2 11396 10556 11396 10556 0 clknet_0_clk
rlabel metal2 6356 11060 6356 11060 0 clknet_1_0__leaf_clk
rlabel metal3 11116 13468 11116 13468 0 clknet_1_1__leaf_clk
rlabel metal3 7140 8428 7140 8428 0 dut6.count\[0\]
rlabel metal2 7784 8316 7784 8316 0 dut6.count\[1\]
rlabel metal2 9968 12012 9968 12012 0 dut6.count\[2\]
rlabel metal2 6748 10696 6748 10696 0 dut6.count\[3\]
rlabel metal3 3178 9604 3178 9604 0 net1
rlabel metal3 3178 11564 3178 11564 0 net10
rlabel metal3 14714 13188 14714 13188 0 net11
rlabel metal2 13468 12768 13468 12768 0 net12
rlabel metal2 13580 8652 13580 8652 0 net13
rlabel metal3 9156 7308 9156 7308 0 net14
rlabel metal2 10164 14056 10164 14056 0 net15
rlabel metal3 18844 10808 18844 10808 0 net16
rlabel metal2 5740 12712 5740 12712 0 net17
rlabel metal3 15960 9688 15960 9688 0 net18
rlabel metal2 14700 9380 14700 9380 0 net19
rlabel metal2 11508 13496 11508 13496 0 net2
rlabel metal2 6524 11732 6524 11732 0 net20
rlabel metal2 9212 13664 9212 13664 0 net21
rlabel metal2 13804 11340 13804 11340 0 net22
rlabel metal2 12628 3178 12628 3178 0 net23
rlabel metal2 10556 2982 10556 2982 0 net24
rlabel metal2 20132 13272 20132 13272 0 net25
rlabel metal2 10108 1015 10108 1015 0 net26
rlabel metal2 11732 13720 11732 13720 0 net3
rlabel metal2 12292 2982 12292 2982 0 net4
rlabel metal3 18844 12376 18844 12376 0 net5
rlabel metal2 18956 10752 18956 10752 0 net6
rlabel metal3 15960 12320 15960 12320 0 net7
rlabel metal2 14980 10752 14980 10752 0 net8
rlabel metal2 2156 13496 2156 13496 0 net9
rlabel metal3 679 9436 679 9436 0 segm[10]
rlabel metal2 11116 19845 11116 19845 0 segm[11]
rlabel metal2 12124 19873 12124 19873 0 segm[12]
rlabel metal2 11452 1099 11452 1099 0 segm[13]
rlabel metal2 20020 12180 20020 12180 0 segm[1]
rlabel metal2 20020 11172 20020 11172 0 segm[2]
rlabel metal2 20020 11900 20020 11900 0 segm[4]
rlabel metal3 20321 10444 20321 10444 0 segm[5]
rlabel metal3 679 13132 679 13132 0 segm[6]
rlabel metal3 679 11452 679 11452 0 segm[7]
rlabel metal2 19964 12936 19964 12936 0 segm[8]
rlabel metal2 20020 12628 20020 12628 0 segm[9]
rlabel metal2 20020 8820 20020 8820 0 sel[0]
rlabel metal2 9436 1211 9436 1211 0 sel[10]
rlabel metal2 9772 19677 9772 19677 0 sel[11]
rlabel metal2 20020 10752 20020 10752 0 sel[1]
rlabel metal3 679 12796 679 12796 0 sel[2]
rlabel metal3 20321 10108 20321 10108 0 sel[3]
rlabel metal2 20020 9548 20020 9548 0 sel[4]
rlabel metal3 679 11788 679 11788 0 sel[5]
rlabel metal2 9100 19873 9100 19873 0 sel[6]
rlabel metal3 20321 11452 20321 11452 0 sel[7]
rlabel metal2 12460 1211 12460 1211 0 sel[8]
rlabel metal2 10444 1099 10444 1099 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
