magic
tech gf180mcuD
magscale 1 10
timestamp 1699642669
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 39790 36370 39842 36382
rect 39790 36306 39842 36318
rect 40238 36258 40290 36270
rect 40238 36194 40290 36206
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 24210 27134 24222 27186
rect 24274 27134 24286 27186
rect 21410 27022 21422 27074
rect 21474 27022 21486 27074
rect 20414 26962 20466 26974
rect 20414 26898 20466 26910
rect 20638 26962 20690 26974
rect 20638 26898 20690 26910
rect 20750 26962 20802 26974
rect 24670 26962 24722 26974
rect 22082 26910 22094 26962
rect 22146 26910 22158 26962
rect 20750 26898 20802 26910
rect 24670 26898 24722 26910
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 25342 26514 25394 26526
rect 25342 26450 25394 26462
rect 17490 26238 17502 26290
rect 17554 26238 17566 26290
rect 21858 26238 21870 26290
rect 21922 26238 21934 26290
rect 16942 26178 16994 26190
rect 18162 26126 18174 26178
rect 18226 26126 18238 26178
rect 20290 26126 20302 26178
rect 20354 26126 20366 26178
rect 22530 26126 22542 26178
rect 22594 26126 22606 26178
rect 24658 26126 24670 26178
rect 24722 26126 24734 26178
rect 16942 26114 16994 26126
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 22766 25730 22818 25742
rect 22766 25666 22818 25678
rect 1934 25618 1986 25630
rect 19518 25618 19570 25630
rect 19058 25566 19070 25618
rect 19122 25566 19134 25618
rect 1934 25554 1986 25566
rect 19518 25554 19570 25566
rect 20414 25618 20466 25630
rect 20414 25554 20466 25566
rect 40014 25618 40066 25630
rect 40014 25554 40066 25566
rect 20078 25506 20130 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 16258 25454 16270 25506
rect 16322 25454 16334 25506
rect 20078 25442 20130 25454
rect 23102 25506 23154 25518
rect 23102 25442 23154 25454
rect 23438 25506 23490 25518
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 23438 25442 23490 25454
rect 22654 25394 22706 25406
rect 16930 25342 16942 25394
rect 16994 25342 17006 25394
rect 22654 25330 22706 25342
rect 23326 25394 23378 25406
rect 23326 25330 23378 25342
rect 23998 25394 24050 25406
rect 23998 25330 24050 25342
rect 24110 25394 24162 25406
rect 24110 25330 24162 25342
rect 19406 25282 19458 25294
rect 19406 25218 19458 25230
rect 19630 25282 19682 25294
rect 19630 25218 19682 25230
rect 22766 25282 22818 25294
rect 22766 25218 22818 25230
rect 23774 25282 23826 25294
rect 23774 25218 23826 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 16158 24946 16210 24958
rect 15362 24894 15374 24946
rect 15426 24894 15438 24946
rect 16158 24882 16210 24894
rect 18286 24946 18338 24958
rect 18286 24882 18338 24894
rect 18622 24946 18674 24958
rect 18622 24882 18674 24894
rect 20526 24946 20578 24958
rect 20526 24882 20578 24894
rect 20190 24834 20242 24846
rect 20190 24770 20242 24782
rect 20302 24834 20354 24846
rect 20302 24770 20354 24782
rect 24446 24834 24498 24846
rect 24446 24770 24498 24782
rect 25342 24834 25394 24846
rect 25342 24770 25394 24782
rect 18174 24722 18226 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 15026 24670 15038 24722
rect 15090 24670 15102 24722
rect 15586 24670 15598 24722
rect 15650 24670 15662 24722
rect 18174 24658 18226 24670
rect 18398 24722 18450 24734
rect 18398 24658 18450 24670
rect 19854 24722 19906 24734
rect 19854 24658 19906 24670
rect 24558 24722 24610 24734
rect 24558 24658 24610 24670
rect 25230 24722 25282 24734
rect 25230 24658 25282 24670
rect 25566 24722 25618 24734
rect 25566 24658 25618 24670
rect 12114 24558 12126 24610
rect 12178 24558 12190 24610
rect 14242 24558 14254 24610
rect 14306 24558 14318 24610
rect 19394 24558 19406 24610
rect 19458 24558 19470 24610
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 24446 24498 24498 24510
rect 24446 24434 24498 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 19182 24162 19234 24174
rect 19182 24098 19234 24110
rect 13582 24050 13634 24062
rect 24658 23998 24670 24050
rect 24722 23998 24734 24050
rect 26786 23998 26798 24050
rect 26850 23998 26862 24050
rect 13582 23986 13634 23998
rect 20638 23938 20690 23950
rect 14466 23886 14478 23938
rect 14530 23886 14542 23938
rect 20066 23886 20078 23938
rect 20130 23886 20142 23938
rect 20638 23874 20690 23886
rect 20750 23938 20802 23950
rect 23874 23886 23886 23938
rect 23938 23886 23950 23938
rect 20750 23874 20802 23886
rect 14814 23826 14866 23838
rect 14814 23762 14866 23774
rect 19406 23826 19458 23838
rect 20290 23774 20302 23826
rect 20354 23774 20366 23826
rect 19406 23762 19458 23774
rect 14702 23714 14754 23726
rect 14702 23650 14754 23662
rect 19294 23714 19346 23726
rect 19294 23650 19346 23662
rect 27246 23714 27298 23726
rect 27246 23650 27298 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 14242 23326 14254 23378
rect 14306 23326 14318 23378
rect 18834 23326 18846 23378
rect 18898 23326 18910 23378
rect 20302 23322 20354 23334
rect 23314 23326 23326 23378
rect 23378 23326 23390 23378
rect 18398 23266 18450 23278
rect 19618 23214 19630 23266
rect 19682 23214 19694 23266
rect 20302 23258 20354 23270
rect 20414 23266 20466 23278
rect 18398 23202 18450 23214
rect 20414 23202 20466 23214
rect 20974 23266 21026 23278
rect 20974 23202 21026 23214
rect 25230 23266 25282 23278
rect 25230 23202 25282 23214
rect 25342 23266 25394 23278
rect 25342 23202 25394 23214
rect 13918 23154 13970 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 13234 23102 13246 23154
rect 13298 23102 13310 23154
rect 13918 23090 13970 23102
rect 14254 23154 14306 23166
rect 18510 23154 18562 23166
rect 14690 23102 14702 23154
rect 14754 23102 14766 23154
rect 14254 23090 14306 23102
rect 18510 23090 18562 23102
rect 19182 23154 19234 23166
rect 20862 23154 20914 23166
rect 19842 23102 19854 23154
rect 19906 23102 19918 23154
rect 19182 23090 19234 23102
rect 20862 23090 20914 23102
rect 22990 23154 23042 23166
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 22990 23090 23042 23102
rect 10322 22990 10334 23042
rect 10386 22990 10398 23042
rect 12450 22990 12462 23042
rect 12514 22990 12526 23042
rect 1934 22930 1986 22942
rect 20414 22930 20466 22942
rect 14466 22878 14478 22930
rect 14530 22878 14542 22930
rect 1934 22866 1986 22878
rect 20414 22866 20466 22878
rect 20974 22930 21026 22942
rect 20974 22866 21026 22878
rect 25342 22930 25394 22942
rect 25342 22866 25394 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 12462 22594 12514 22606
rect 12462 22530 12514 22542
rect 17950 22594 18002 22606
rect 17950 22530 18002 22542
rect 21310 22594 21362 22606
rect 21310 22530 21362 22542
rect 21646 22594 21698 22606
rect 21646 22530 21698 22542
rect 17390 22482 17442 22494
rect 16930 22430 16942 22482
rect 16994 22430 17006 22482
rect 26338 22430 26350 22482
rect 26402 22430 26414 22482
rect 17390 22418 17442 22430
rect 20190 22370 20242 22382
rect 14130 22318 14142 22370
rect 14194 22318 14206 22370
rect 20190 22306 20242 22318
rect 22206 22370 22258 22382
rect 26798 22370 26850 22382
rect 23538 22318 23550 22370
rect 23602 22318 23614 22370
rect 22206 22306 22258 22318
rect 26798 22306 26850 22318
rect 12574 22258 12626 22270
rect 12574 22194 12626 22206
rect 12798 22258 12850 22270
rect 12798 22194 12850 22206
rect 13582 22258 13634 22270
rect 17838 22258 17890 22270
rect 14802 22206 14814 22258
rect 14866 22206 14878 22258
rect 13582 22194 13634 22206
rect 17838 22194 17890 22206
rect 17950 22258 18002 22270
rect 17950 22194 18002 22206
rect 18510 22258 18562 22270
rect 18510 22194 18562 22206
rect 22094 22258 22146 22270
rect 22094 22194 22146 22206
rect 22766 22258 22818 22270
rect 24210 22206 24222 22258
rect 24274 22206 24286 22258
rect 22766 22194 22818 22206
rect 13694 22146 13746 22158
rect 13694 22082 13746 22094
rect 18398 22146 18450 22158
rect 18398 22082 18450 22094
rect 19518 22146 19570 22158
rect 21534 22146 21586 22158
rect 19842 22094 19854 22146
rect 19906 22094 19918 22146
rect 20514 22094 20526 22146
rect 20578 22094 20590 22146
rect 19518 22082 19570 22094
rect 21534 22082 21586 22094
rect 21870 22146 21922 22158
rect 23090 22094 23102 22146
rect 23154 22094 23166 22146
rect 21870 22082 21922 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 13694 21810 13746 21822
rect 13694 21746 13746 21758
rect 13806 21810 13858 21822
rect 13806 21746 13858 21758
rect 14030 21810 14082 21822
rect 14030 21746 14082 21758
rect 14590 21810 14642 21822
rect 14590 21746 14642 21758
rect 23438 21810 23490 21822
rect 23438 21746 23490 21758
rect 23998 21810 24050 21822
rect 23998 21746 24050 21758
rect 24110 21810 24162 21822
rect 24110 21746 24162 21758
rect 24334 21810 24386 21822
rect 24334 21746 24386 21758
rect 25790 21810 25842 21822
rect 25790 21746 25842 21758
rect 13470 21698 13522 21710
rect 23326 21698 23378 21710
rect 19842 21646 19854 21698
rect 19906 21646 19918 21698
rect 21074 21646 21086 21698
rect 21138 21646 21150 21698
rect 21970 21646 21982 21698
rect 22034 21646 22046 21698
rect 13470 21634 13522 21646
rect 23326 21634 23378 21646
rect 26798 21698 26850 21710
rect 26798 21634 26850 21646
rect 13918 21586 13970 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 13122 21534 13134 21586
rect 13186 21534 13198 21586
rect 13918 21522 13970 21534
rect 17502 21586 17554 21598
rect 17502 21522 17554 21534
rect 18510 21586 18562 21598
rect 22766 21586 22818 21598
rect 23886 21586 23938 21598
rect 20290 21534 20302 21586
rect 20354 21534 20366 21586
rect 22194 21534 22206 21586
rect 22258 21534 22270 21586
rect 23090 21534 23102 21586
rect 23154 21534 23166 21586
rect 18510 21522 18562 21534
rect 22766 21522 22818 21534
rect 23886 21522 23938 21534
rect 25566 21586 25618 21598
rect 25566 21522 25618 21534
rect 26238 21586 26290 21598
rect 26238 21522 26290 21534
rect 26574 21586 26626 21598
rect 26574 21522 26626 21534
rect 26910 21586 26962 21598
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 26910 21522 26962 21534
rect 25678 21474 25730 21486
rect 10210 21422 10222 21474
rect 10274 21422 10286 21474
rect 12338 21422 12350 21474
rect 12402 21422 12414 21474
rect 21298 21422 21310 21474
rect 21362 21422 21374 21474
rect 25678 21410 25730 21422
rect 1934 21362 1986 21374
rect 1934 21298 1986 21310
rect 17726 21362 17778 21374
rect 40014 21362 40066 21374
rect 18050 21310 18062 21362
rect 18114 21310 18126 21362
rect 17726 21298 17778 21310
rect 40014 21298 40066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 12574 21026 12626 21038
rect 12574 20962 12626 20974
rect 12910 21026 12962 21038
rect 12910 20962 12962 20974
rect 17826 20862 17838 20914
rect 17890 20862 17902 20914
rect 18610 20862 18622 20914
rect 18674 20862 18686 20914
rect 25218 20862 25230 20914
rect 25282 20862 25294 20914
rect 13694 20802 13746 20814
rect 13458 20750 13470 20802
rect 13522 20750 13534 20802
rect 13694 20738 13746 20750
rect 13918 20802 13970 20814
rect 18174 20802 18226 20814
rect 20526 20802 20578 20814
rect 16370 20750 16382 20802
rect 16434 20750 16446 20802
rect 17042 20750 17054 20802
rect 17106 20750 17118 20802
rect 18946 20750 18958 20802
rect 19010 20750 19022 20802
rect 19506 20750 19518 20802
rect 19570 20750 19582 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 13918 20738 13970 20750
rect 18174 20738 18226 20750
rect 20526 20738 20578 20750
rect 20862 20802 20914 20814
rect 20862 20738 20914 20750
rect 21646 20802 21698 20814
rect 22306 20750 22318 20802
rect 22370 20750 22382 20802
rect 21646 20738 21698 20750
rect 16606 20690 16658 20702
rect 17614 20690 17666 20702
rect 20638 20690 20690 20702
rect 17266 20638 17278 20690
rect 17330 20638 17342 20690
rect 18834 20638 18846 20690
rect 18898 20638 18910 20690
rect 16606 20626 16658 20638
rect 17614 20626 17666 20638
rect 20638 20626 20690 20638
rect 12686 20578 12738 20590
rect 12686 20514 12738 20526
rect 13806 20578 13858 20590
rect 13806 20514 13858 20526
rect 14030 20578 14082 20590
rect 14030 20514 14082 20526
rect 17838 20578 17890 20590
rect 19842 20526 19854 20578
rect 19906 20526 19918 20578
rect 21970 20526 21982 20578
rect 22034 20526 22046 20578
rect 17838 20514 17890 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 18174 20242 18226 20254
rect 18174 20178 18226 20190
rect 16606 20130 16658 20142
rect 15586 20078 15598 20130
rect 15650 20078 15662 20130
rect 16606 20066 16658 20078
rect 17390 20130 17442 20142
rect 17714 20078 17726 20130
rect 17778 20078 17790 20130
rect 22306 20078 22318 20130
rect 22370 20078 22382 20130
rect 26338 20078 26350 20130
rect 26402 20078 26414 20130
rect 17390 20066 17442 20078
rect 15810 19966 15822 20018
rect 15874 19966 15886 20018
rect 18722 19966 18734 20018
rect 18786 19966 18798 20018
rect 25554 19966 25566 20018
rect 25618 19966 25630 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 18398 19906 18450 19918
rect 28926 19906 28978 19918
rect 18050 19854 18062 19906
rect 18114 19854 18126 19906
rect 28466 19854 28478 19906
rect 28530 19854 28542 19906
rect 18398 19842 18450 19854
rect 28926 19842 28978 19854
rect 16494 19794 16546 19806
rect 16494 19730 16546 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 24110 19458 24162 19470
rect 22082 19406 22094 19458
rect 22146 19406 22158 19458
rect 24110 19394 24162 19406
rect 14254 19346 14306 19358
rect 14690 19294 14702 19346
rect 14754 19294 14766 19346
rect 24434 19294 24446 19346
rect 24498 19294 24510 19346
rect 26002 19294 26014 19346
rect 26066 19294 26078 19346
rect 28130 19294 28142 19346
rect 28194 19294 28206 19346
rect 14254 19282 14306 19294
rect 14030 19234 14082 19246
rect 21422 19234 21474 19246
rect 22766 19234 22818 19246
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 14030 19170 14082 19182
rect 21422 19170 21474 19182
rect 22766 19170 22818 19182
rect 23102 19234 23154 19246
rect 23102 19170 23154 19182
rect 23438 19234 23490 19246
rect 23438 19170 23490 19182
rect 23886 19234 23938 19246
rect 23886 19170 23938 19182
rect 24558 19234 24610 19246
rect 25218 19182 25230 19234
rect 25282 19182 25294 19234
rect 24558 19170 24610 19182
rect 12910 19122 12962 19134
rect 12910 19058 12962 19070
rect 14702 19122 14754 19134
rect 14702 19058 14754 19070
rect 14926 19122 14978 19134
rect 24670 19122 24722 19134
rect 15474 19070 15486 19122
rect 15538 19070 15550 19122
rect 14926 19058 14978 19070
rect 24670 19058 24722 19070
rect 12574 19010 12626 19022
rect 22990 19010 23042 19022
rect 13682 18958 13694 19010
rect 13746 18958 13758 19010
rect 12574 18946 12626 18958
rect 22990 18946 23042 18958
rect 28590 19010 28642 19022
rect 28590 18946 28642 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 17950 18674 18002 18686
rect 17950 18610 18002 18622
rect 18174 18674 18226 18686
rect 18174 18610 18226 18622
rect 26574 18674 26626 18686
rect 26574 18610 26626 18622
rect 18286 18562 18338 18574
rect 25902 18562 25954 18574
rect 12226 18510 12238 18562
rect 12290 18510 12302 18562
rect 16258 18510 16270 18562
rect 16322 18510 16334 18562
rect 18498 18510 18510 18562
rect 18562 18510 18574 18562
rect 19394 18510 19406 18562
rect 19458 18510 19470 18562
rect 18286 18498 18338 18510
rect 25902 18498 25954 18510
rect 26686 18562 26738 18574
rect 26686 18498 26738 18510
rect 27022 18562 27074 18574
rect 27022 18498 27074 18510
rect 27134 18562 27186 18574
rect 27134 18498 27186 18510
rect 14814 18450 14866 18462
rect 17726 18450 17778 18462
rect 20638 18450 20690 18462
rect 11554 18398 11566 18450
rect 11618 18398 11630 18450
rect 16034 18398 16046 18450
rect 16098 18398 16110 18450
rect 19058 18398 19070 18450
rect 19122 18398 19134 18450
rect 19954 18398 19966 18450
rect 20018 18398 20030 18450
rect 14814 18386 14866 18398
rect 17726 18386 17778 18398
rect 20638 18386 20690 18398
rect 25342 18450 25394 18462
rect 25342 18386 25394 18398
rect 26350 18450 26402 18462
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 26350 18386 26402 18398
rect 18062 18338 18114 18350
rect 20974 18338 21026 18350
rect 14354 18286 14366 18338
rect 14418 18286 14430 18338
rect 19506 18286 19518 18338
rect 19570 18286 19582 18338
rect 25778 18286 25790 18338
rect 25842 18286 25854 18338
rect 18062 18274 18114 18286
rect 20974 18274 21026 18286
rect 20526 18226 20578 18238
rect 20526 18162 20578 18174
rect 20862 18226 20914 18238
rect 20862 18162 20914 18174
rect 25566 18226 25618 18238
rect 25566 18162 25618 18174
rect 26126 18226 26178 18238
rect 26126 18162 26178 18174
rect 27134 18226 27186 18238
rect 27134 18162 27186 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 21422 17890 21474 17902
rect 21422 17826 21474 17838
rect 21646 17890 21698 17902
rect 21646 17826 21698 17838
rect 22094 17890 22146 17902
rect 22094 17826 22146 17838
rect 1934 17778 1986 17790
rect 16158 17778 16210 17790
rect 15698 17726 15710 17778
rect 15762 17726 15774 17778
rect 25554 17726 25566 17778
rect 25618 17726 25630 17778
rect 27682 17726 27694 17778
rect 27746 17726 27758 17778
rect 1934 17714 1986 17726
rect 16158 17714 16210 17726
rect 15598 17666 15650 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 15138 17614 15150 17666
rect 15202 17614 15214 17666
rect 15598 17602 15650 17614
rect 18622 17666 18674 17678
rect 20190 17666 20242 17678
rect 19842 17614 19854 17666
rect 19906 17614 19918 17666
rect 18622 17602 18674 17614
rect 20190 17602 20242 17614
rect 20638 17666 20690 17678
rect 20638 17602 20690 17614
rect 21982 17666 22034 17678
rect 21982 17602 22034 17614
rect 22430 17666 22482 17678
rect 22430 17602 22482 17614
rect 22766 17666 22818 17678
rect 22766 17602 22818 17614
rect 22990 17666 23042 17678
rect 24770 17614 24782 17666
rect 24834 17614 24846 17666
rect 22990 17602 23042 17614
rect 15374 17554 15426 17566
rect 15374 17490 15426 17502
rect 18398 17554 18450 17566
rect 18398 17490 18450 17502
rect 18846 17554 18898 17566
rect 22206 17554 22258 17566
rect 20402 17502 20414 17554
rect 20466 17502 20478 17554
rect 18846 17490 18898 17502
rect 22206 17490 22258 17502
rect 15710 17442 15762 17454
rect 15710 17378 15762 17390
rect 16270 17442 16322 17454
rect 16270 17378 16322 17390
rect 16382 17442 16434 17454
rect 16382 17378 16434 17390
rect 18734 17442 18786 17454
rect 18734 17378 18786 17390
rect 19854 17442 19906 17454
rect 19854 17378 19906 17390
rect 22766 17442 22818 17454
rect 22766 17378 22818 17390
rect 28142 17442 28194 17454
rect 28142 17378 28194 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 17278 17106 17330 17118
rect 17278 17042 17330 17054
rect 17502 17106 17554 17118
rect 17502 17042 17554 17054
rect 20190 17106 20242 17118
rect 20190 17042 20242 17054
rect 22094 17106 22146 17118
rect 22094 17042 22146 17054
rect 22318 17106 22370 17118
rect 22318 17042 22370 17054
rect 16606 16994 16658 17006
rect 14578 16942 14590 16994
rect 14642 16942 14654 16994
rect 16606 16930 16658 16942
rect 17614 16994 17666 17006
rect 17614 16930 17666 16942
rect 20078 16994 20130 17006
rect 20078 16930 20130 16942
rect 21982 16994 22034 17006
rect 25554 16942 25566 16994
rect 25618 16942 25630 16994
rect 21982 16930 22034 16942
rect 15822 16882 15874 16894
rect 15362 16830 15374 16882
rect 15426 16830 15438 16882
rect 15822 16818 15874 16830
rect 16158 16882 16210 16894
rect 16158 16818 16210 16830
rect 16494 16882 16546 16894
rect 16494 16818 16546 16830
rect 16830 16882 16882 16894
rect 16830 16818 16882 16830
rect 20302 16882 20354 16894
rect 20302 16818 20354 16830
rect 20750 16882 20802 16894
rect 25330 16830 25342 16882
rect 25394 16830 25406 16882
rect 20750 16818 20802 16830
rect 20526 16770 20578 16782
rect 12450 16718 12462 16770
rect 12514 16718 12526 16770
rect 20526 16706 20578 16718
rect 20974 16770 21026 16782
rect 20974 16706 21026 16718
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 17502 16210 17554 16222
rect 26350 16210 26402 16222
rect 14690 16158 14702 16210
rect 14754 16158 14766 16210
rect 16818 16158 16830 16210
rect 16882 16158 16894 16210
rect 18610 16158 18622 16210
rect 18674 16158 18686 16210
rect 20738 16158 20750 16210
rect 20802 16158 20814 16210
rect 23538 16158 23550 16210
rect 23602 16158 23614 16210
rect 17502 16146 17554 16158
rect 26350 16146 26402 16158
rect 14018 16046 14030 16098
rect 14082 16046 14094 16098
rect 17826 16046 17838 16098
rect 17890 16046 17902 16098
rect 22866 16046 22878 16098
rect 22930 16046 22942 16098
rect 25778 15822 25790 15874
rect 25842 15822 25854 15874
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 17502 15538 17554 15550
rect 21310 15538 21362 15550
rect 20962 15486 20974 15538
rect 21026 15486 21038 15538
rect 17502 15474 17554 15486
rect 21310 15474 21362 15486
rect 20078 15426 20130 15438
rect 20078 15362 20130 15374
rect 20638 15426 20690 15438
rect 25554 15374 25566 15426
rect 25618 15374 25630 15426
rect 20638 15362 20690 15374
rect 20414 15314 20466 15326
rect 25330 15262 25342 15314
rect 25394 15262 25406 15314
rect 20414 15250 20466 15262
rect 20190 15202 20242 15214
rect 20190 15138 20242 15150
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19518 14754 19570 14766
rect 19518 14690 19570 14702
rect 21422 14754 21474 14766
rect 21422 14690 21474 14702
rect 21646 14754 21698 14766
rect 21646 14690 21698 14702
rect 17950 14642 18002 14654
rect 17950 14578 18002 14590
rect 22318 14642 22370 14654
rect 22318 14578 22370 14590
rect 16146 14478 16158 14530
rect 16210 14478 16222 14530
rect 19170 14478 19182 14530
rect 19234 14478 19246 14530
rect 21858 14478 21870 14530
rect 21922 14478 21934 14530
rect 22530 14478 22542 14530
rect 22594 14478 22606 14530
rect 16494 14418 16546 14430
rect 16494 14354 16546 14366
rect 22206 14418 22258 14430
rect 22206 14354 22258 14366
rect 16382 14306 16434 14318
rect 16382 14242 16434 14254
rect 17166 14306 17218 14318
rect 19406 14306 19458 14318
rect 17490 14254 17502 14306
rect 17554 14254 17566 14306
rect 17166 14242 17218 14254
rect 19406 14242 19458 14254
rect 21758 14306 21810 14318
rect 21758 14242 21810 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 24110 13970 24162 13982
rect 24110 13906 24162 13918
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 18274 13806 18286 13858
rect 18338 13806 18350 13858
rect 21522 13806 21534 13858
rect 21586 13806 21598 13858
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 17602 13694 17614 13746
rect 17666 13694 17678 13746
rect 20850 13694 20862 13746
rect 20914 13694 20926 13746
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 20402 13582 20414 13634
rect 20466 13582 20478 13634
rect 23650 13582 23662 13634
rect 23714 13582 23726 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 17390 13186 17442 13198
rect 17390 13122 17442 13134
rect 17950 13074 18002 13086
rect 17154 13022 17166 13074
rect 17218 13022 17230 13074
rect 17950 13010 18002 13022
rect 22978 12910 22990 12962
rect 23042 12910 23054 12962
rect 17166 12850 17218 12862
rect 17166 12786 17218 12798
rect 23202 12686 23214 12738
rect 23266 12686 23278 12738
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 20402 5854 20414 5906
rect 20466 5854 20478 5906
rect 21422 5682 21474 5694
rect 21422 5618 21474 5630
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 18062 5234 18114 5246
rect 18062 5170 18114 5182
rect 24782 5234 24834 5246
rect 24782 5170 24834 5182
rect 17042 5070 17054 5122
rect 17106 5070 17118 5122
rect 23762 5070 23774 5122
rect 23826 5070 23838 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 17266 4398 17278 4450
rect 17330 4447 17342 4450
rect 17602 4447 17614 4450
rect 17330 4401 17614 4447
rect 17330 4398 17342 4401
rect 17602 4398 17614 4401
rect 17666 4398 17678 4450
rect 17714 4286 17726 4338
rect 17778 4286 17790 4338
rect 21074 4286 21086 4338
rect 21138 4286 21150 4338
rect 25554 4286 25566 4338
rect 25618 4286 25630 4338
rect 18734 4114 18786 4126
rect 18734 4050 18786 4062
rect 22094 4114 22146 4126
rect 22094 4050 22146 4062
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 23650 3502 23662 3554
rect 23714 3502 23726 3554
rect 24994 3502 25006 3554
rect 25058 3502 25070 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 22194 3390 22206 3442
rect 22258 3390 22270 3442
rect 21086 3330 21138 3342
rect 21086 3266 21138 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 25566 38222 25618 38274
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 26238 37438 26290 37490
rect 25230 37214 25282 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 1710 36318 1762 36370
rect 39790 36318 39842 36370
rect 40238 36206 40290 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 24222 27134 24274 27186
rect 21422 27022 21474 27074
rect 20414 26910 20466 26962
rect 20638 26910 20690 26962
rect 20750 26910 20802 26962
rect 22094 26910 22146 26962
rect 24670 26910 24722 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 25342 26462 25394 26514
rect 17502 26238 17554 26290
rect 21870 26238 21922 26290
rect 16942 26126 16994 26178
rect 18174 26126 18226 26178
rect 20302 26126 20354 26178
rect 22542 26126 22594 26178
rect 24670 26126 24722 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 22766 25678 22818 25730
rect 1934 25566 1986 25618
rect 19070 25566 19122 25618
rect 19518 25566 19570 25618
rect 20414 25566 20466 25618
rect 40014 25566 40066 25618
rect 4286 25454 4338 25506
rect 16270 25454 16322 25506
rect 20078 25454 20130 25506
rect 23102 25454 23154 25506
rect 23438 25454 23490 25506
rect 37662 25454 37714 25506
rect 16942 25342 16994 25394
rect 22654 25342 22706 25394
rect 23326 25342 23378 25394
rect 23998 25342 24050 25394
rect 24110 25342 24162 25394
rect 19406 25230 19458 25282
rect 19630 25230 19682 25282
rect 22766 25230 22818 25282
rect 23774 25230 23826 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 15374 24894 15426 24946
rect 16158 24894 16210 24946
rect 18286 24894 18338 24946
rect 18622 24894 18674 24946
rect 20526 24894 20578 24946
rect 20190 24782 20242 24834
rect 20302 24782 20354 24834
rect 24446 24782 24498 24834
rect 25342 24782 25394 24834
rect 4286 24670 4338 24722
rect 15038 24670 15090 24722
rect 15598 24670 15650 24722
rect 18174 24670 18226 24722
rect 18398 24670 18450 24722
rect 19854 24670 19906 24722
rect 24558 24670 24610 24722
rect 25230 24670 25282 24722
rect 25566 24670 25618 24722
rect 12126 24558 12178 24610
rect 14254 24558 14306 24610
rect 19406 24558 19458 24610
rect 1934 24446 1986 24498
rect 24446 24446 24498 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 19182 24110 19234 24162
rect 13582 23998 13634 24050
rect 24670 23998 24722 24050
rect 26798 23998 26850 24050
rect 14478 23886 14530 23938
rect 20078 23886 20130 23938
rect 20638 23886 20690 23938
rect 20750 23886 20802 23938
rect 23886 23886 23938 23938
rect 14814 23774 14866 23826
rect 19406 23774 19458 23826
rect 20302 23774 20354 23826
rect 14702 23662 14754 23714
rect 19294 23662 19346 23714
rect 27246 23662 27298 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 14254 23326 14306 23378
rect 18846 23326 18898 23378
rect 23326 23326 23378 23378
rect 20302 23270 20354 23322
rect 18398 23214 18450 23266
rect 19630 23214 19682 23266
rect 20414 23214 20466 23266
rect 20974 23214 21026 23266
rect 25230 23214 25282 23266
rect 25342 23214 25394 23266
rect 4286 23102 4338 23154
rect 13246 23102 13298 23154
rect 13918 23102 13970 23154
rect 14254 23102 14306 23154
rect 14702 23102 14754 23154
rect 18510 23102 18562 23154
rect 19182 23102 19234 23154
rect 19854 23102 19906 23154
rect 20862 23102 20914 23154
rect 22990 23102 23042 23154
rect 37662 23102 37714 23154
rect 10334 22990 10386 23042
rect 12462 22990 12514 23042
rect 1934 22878 1986 22930
rect 14478 22878 14530 22930
rect 20414 22878 20466 22930
rect 20974 22878 21026 22930
rect 25342 22878 25394 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 12462 22542 12514 22594
rect 17950 22542 18002 22594
rect 21310 22542 21362 22594
rect 21646 22542 21698 22594
rect 16942 22430 16994 22482
rect 17390 22430 17442 22482
rect 26350 22430 26402 22482
rect 14142 22318 14194 22370
rect 20190 22318 20242 22370
rect 22206 22318 22258 22370
rect 23550 22318 23602 22370
rect 26798 22318 26850 22370
rect 12574 22206 12626 22258
rect 12798 22206 12850 22258
rect 13582 22206 13634 22258
rect 14814 22206 14866 22258
rect 17838 22206 17890 22258
rect 17950 22206 18002 22258
rect 18510 22206 18562 22258
rect 22094 22206 22146 22258
rect 22766 22206 22818 22258
rect 24222 22206 24274 22258
rect 13694 22094 13746 22146
rect 18398 22094 18450 22146
rect 19518 22094 19570 22146
rect 19854 22094 19906 22146
rect 20526 22094 20578 22146
rect 21534 22094 21586 22146
rect 21870 22094 21922 22146
rect 23102 22094 23154 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 13694 21758 13746 21810
rect 13806 21758 13858 21810
rect 14030 21758 14082 21810
rect 14590 21758 14642 21810
rect 23438 21758 23490 21810
rect 23998 21758 24050 21810
rect 24110 21758 24162 21810
rect 24334 21758 24386 21810
rect 25790 21758 25842 21810
rect 13470 21646 13522 21698
rect 19854 21646 19906 21698
rect 21086 21646 21138 21698
rect 21982 21646 22034 21698
rect 23326 21646 23378 21698
rect 26798 21646 26850 21698
rect 4286 21534 4338 21586
rect 13134 21534 13186 21586
rect 13918 21534 13970 21586
rect 17502 21534 17554 21586
rect 18510 21534 18562 21586
rect 20302 21534 20354 21586
rect 22206 21534 22258 21586
rect 22766 21534 22818 21586
rect 23102 21534 23154 21586
rect 23886 21534 23938 21586
rect 25566 21534 25618 21586
rect 26238 21534 26290 21586
rect 26574 21534 26626 21586
rect 26910 21534 26962 21586
rect 37662 21534 37714 21586
rect 10222 21422 10274 21474
rect 12350 21422 12402 21474
rect 21310 21422 21362 21474
rect 25678 21422 25730 21474
rect 1934 21310 1986 21362
rect 17726 21310 17778 21362
rect 18062 21310 18114 21362
rect 40014 21310 40066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 12574 20974 12626 21026
rect 12910 20974 12962 21026
rect 17838 20862 17890 20914
rect 18622 20862 18674 20914
rect 25230 20862 25282 20914
rect 13470 20750 13522 20802
rect 13694 20750 13746 20802
rect 13918 20750 13970 20802
rect 16382 20750 16434 20802
rect 17054 20750 17106 20802
rect 18174 20750 18226 20802
rect 18958 20750 19010 20802
rect 19518 20750 19570 20802
rect 20078 20750 20130 20802
rect 20526 20750 20578 20802
rect 20862 20750 20914 20802
rect 21646 20750 21698 20802
rect 22318 20750 22370 20802
rect 16606 20638 16658 20690
rect 17278 20638 17330 20690
rect 17614 20638 17666 20690
rect 18846 20638 18898 20690
rect 20638 20638 20690 20690
rect 12686 20526 12738 20578
rect 13806 20526 13858 20578
rect 14030 20526 14082 20578
rect 17838 20526 17890 20578
rect 19854 20526 19906 20578
rect 21982 20526 22034 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 18174 20190 18226 20242
rect 15598 20078 15650 20130
rect 16606 20078 16658 20130
rect 17390 20078 17442 20130
rect 17726 20078 17778 20130
rect 22318 20078 22370 20130
rect 26350 20078 26402 20130
rect 15822 19966 15874 20018
rect 18734 19966 18786 20018
rect 25566 19966 25618 20018
rect 37662 19966 37714 20018
rect 18062 19854 18114 19906
rect 18398 19854 18450 19906
rect 28478 19854 28530 19906
rect 28926 19854 28978 19906
rect 16494 19742 16546 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 22094 19406 22146 19458
rect 24110 19406 24162 19458
rect 14254 19294 14306 19346
rect 14702 19294 14754 19346
rect 24446 19294 24498 19346
rect 26014 19294 26066 19346
rect 28142 19294 28194 19346
rect 14030 19182 14082 19234
rect 20078 19182 20130 19234
rect 21422 19182 21474 19234
rect 21758 19182 21810 19234
rect 22766 19182 22818 19234
rect 23102 19182 23154 19234
rect 23438 19182 23490 19234
rect 23886 19182 23938 19234
rect 24558 19182 24610 19234
rect 25230 19182 25282 19234
rect 12910 19070 12962 19122
rect 14702 19070 14754 19122
rect 14926 19070 14978 19122
rect 15486 19070 15538 19122
rect 24670 19070 24722 19122
rect 12574 18958 12626 19010
rect 13694 18958 13746 19010
rect 22990 18958 23042 19010
rect 28590 18958 28642 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 17950 18622 18002 18674
rect 18174 18622 18226 18674
rect 26574 18622 26626 18674
rect 12238 18510 12290 18562
rect 16270 18510 16322 18562
rect 18286 18510 18338 18562
rect 18510 18510 18562 18562
rect 19406 18510 19458 18562
rect 25902 18510 25954 18562
rect 26686 18510 26738 18562
rect 27022 18510 27074 18562
rect 27134 18510 27186 18562
rect 11566 18398 11618 18450
rect 14814 18398 14866 18450
rect 16046 18398 16098 18450
rect 17726 18398 17778 18450
rect 19070 18398 19122 18450
rect 19966 18398 20018 18450
rect 20638 18398 20690 18450
rect 25342 18398 25394 18450
rect 26350 18398 26402 18450
rect 37662 18398 37714 18450
rect 14366 18286 14418 18338
rect 18062 18286 18114 18338
rect 19518 18286 19570 18338
rect 20974 18286 21026 18338
rect 25790 18286 25842 18338
rect 20526 18174 20578 18226
rect 20862 18174 20914 18226
rect 25566 18174 25618 18226
rect 26126 18174 26178 18226
rect 27134 18174 27186 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 21422 17838 21474 17890
rect 21646 17838 21698 17890
rect 22094 17838 22146 17890
rect 1934 17726 1986 17778
rect 15710 17726 15762 17778
rect 16158 17726 16210 17778
rect 25566 17726 25618 17778
rect 27694 17726 27746 17778
rect 4286 17614 4338 17666
rect 15150 17614 15202 17666
rect 15598 17614 15650 17666
rect 18622 17614 18674 17666
rect 19854 17614 19906 17666
rect 20190 17614 20242 17666
rect 20638 17614 20690 17666
rect 21982 17614 22034 17666
rect 22430 17614 22482 17666
rect 22766 17614 22818 17666
rect 22990 17614 23042 17666
rect 24782 17614 24834 17666
rect 15374 17502 15426 17554
rect 18398 17502 18450 17554
rect 18846 17502 18898 17554
rect 20414 17502 20466 17554
rect 22206 17502 22258 17554
rect 15710 17390 15762 17442
rect 16270 17390 16322 17442
rect 16382 17390 16434 17442
rect 18734 17390 18786 17442
rect 19854 17390 19906 17442
rect 22766 17390 22818 17442
rect 28142 17390 28194 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17278 17054 17330 17106
rect 17502 17054 17554 17106
rect 20190 17054 20242 17106
rect 22094 17054 22146 17106
rect 22318 17054 22370 17106
rect 14590 16942 14642 16994
rect 16606 16942 16658 16994
rect 17614 16942 17666 16994
rect 20078 16942 20130 16994
rect 21982 16942 22034 16994
rect 25566 16942 25618 16994
rect 15374 16830 15426 16882
rect 15822 16830 15874 16882
rect 16158 16830 16210 16882
rect 16494 16830 16546 16882
rect 16830 16830 16882 16882
rect 20302 16830 20354 16882
rect 20750 16830 20802 16882
rect 25342 16830 25394 16882
rect 12462 16718 12514 16770
rect 20526 16718 20578 16770
rect 20974 16718 21026 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 14702 16158 14754 16210
rect 16830 16158 16882 16210
rect 17502 16158 17554 16210
rect 18622 16158 18674 16210
rect 20750 16158 20802 16210
rect 23550 16158 23602 16210
rect 26350 16158 26402 16210
rect 14030 16046 14082 16098
rect 17838 16046 17890 16098
rect 22878 16046 22930 16098
rect 25790 15822 25842 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 17502 15486 17554 15538
rect 20974 15486 21026 15538
rect 21310 15486 21362 15538
rect 20078 15374 20130 15426
rect 20638 15374 20690 15426
rect 25566 15374 25618 15426
rect 20414 15262 20466 15314
rect 25342 15262 25394 15314
rect 20190 15150 20242 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19518 14702 19570 14754
rect 21422 14702 21474 14754
rect 21646 14702 21698 14754
rect 17950 14590 18002 14642
rect 22318 14590 22370 14642
rect 16158 14478 16210 14530
rect 19182 14478 19234 14530
rect 21870 14478 21922 14530
rect 22542 14478 22594 14530
rect 16494 14366 16546 14418
rect 22206 14366 22258 14418
rect 16382 14254 16434 14306
rect 17166 14254 17218 14306
rect 17502 14254 17554 14306
rect 19406 14254 19458 14306
rect 21758 14254 21810 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 24110 13918 24162 13970
rect 14702 13806 14754 13858
rect 18286 13806 18338 13858
rect 21534 13806 21586 13858
rect 14030 13694 14082 13746
rect 17614 13694 17666 13746
rect 20862 13694 20914 13746
rect 16830 13582 16882 13634
rect 20414 13582 20466 13634
rect 23662 13582 23714 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17390 13134 17442 13186
rect 17166 13022 17218 13074
rect 17950 13022 18002 13074
rect 22990 12910 23042 12962
rect 17166 12798 17218 12850
rect 23214 12686 23266 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 20414 5854 20466 5906
rect 21422 5630 21474 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 18062 5182 18114 5234
rect 24782 5182 24834 5234
rect 17054 5070 17106 5122
rect 23774 5070 23826 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 17278 4398 17330 4450
rect 17614 4398 17666 4450
rect 17726 4286 17778 4338
rect 21086 4286 21138 4338
rect 25566 4286 25618 4338
rect 18734 4062 18786 4114
rect 22094 4062 22146 4114
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 25566 3614 25618 3666
rect 29374 3614 29426 3666
rect 17614 3502 17666 3554
rect 23662 3502 23714 3554
rect 25006 3502 25058 3554
rect 28590 3502 28642 3554
rect 22206 3390 22258 3442
rect 21086 3278 21138 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 22848 41200 22960 42000
rect 24864 41200 24976 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1708 36372 1764 36382
rect 1708 36278 1764 36316
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 24556 31948 24612 37998
rect 24892 37492 24948 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 24892 37426 24948 37436
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 24220 31892 24612 31948
rect 25228 37266 25284 37278
rect 25228 37214 25230 37266
rect 25282 37214 25284 37266
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 24220 27186 24276 31892
rect 24220 27134 24222 27186
rect 24274 27134 24276 27186
rect 21420 27076 21476 27086
rect 21420 27074 21812 27076
rect 21420 27022 21422 27074
rect 21474 27022 21812 27074
rect 21420 27020 21812 27022
rect 21420 27010 21476 27020
rect 20412 26964 20468 26974
rect 20412 26870 20468 26908
rect 20636 26962 20692 26974
rect 20636 26910 20638 26962
rect 20690 26910 20692 26962
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20636 26404 20692 26910
rect 20076 26348 20692 26404
rect 4172 26292 4228 26302
rect 1932 25618 1988 25630
rect 1932 25566 1934 25618
rect 1986 25566 1988 25618
rect 1932 24948 1988 25566
rect 1932 24882 1988 24892
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 21362 1988 21374
rect 1932 21310 1934 21362
rect 1986 21310 1988 21362
rect 1932 20916 1988 21310
rect 1932 20850 1988 20860
rect 4172 19348 4228 26236
rect 17500 26290 17556 26302
rect 17500 26238 17502 26290
rect 17554 26238 17556 26290
rect 16940 26180 16996 26190
rect 17500 26180 17556 26238
rect 16940 26178 17556 26180
rect 16940 26126 16942 26178
rect 16994 26126 17556 26178
rect 16940 26124 17556 26126
rect 16940 26114 16996 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 16268 25620 16324 25630
rect 17500 25620 17556 26124
rect 18172 26180 18228 26190
rect 18172 26086 18228 26124
rect 19516 26180 19572 26190
rect 4284 25508 4340 25518
rect 4284 25414 4340 25452
rect 15372 25508 15428 25518
rect 16268 25508 16324 25564
rect 13580 24948 13636 24958
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 12124 24724 12180 24734
rect 12124 24610 12180 24668
rect 12124 24558 12126 24610
rect 12178 24558 12180 24610
rect 12124 24546 12180 24558
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 13580 24052 13636 24892
rect 15036 24948 15092 24958
rect 14476 24724 14532 24734
rect 13468 24050 13636 24052
rect 13468 23998 13582 24050
rect 13634 23998 13636 24050
rect 13468 23996 13636 23998
rect 4284 23156 4340 23166
rect 13244 23156 13300 23166
rect 13468 23156 13524 23996
rect 13580 23986 13636 23996
rect 14252 24610 14308 24622
rect 14252 24558 14254 24610
rect 14306 24558 14308 24610
rect 14140 23604 14196 23614
rect 14028 23548 14140 23604
rect 13916 23156 13972 23166
rect 4284 23062 4340 23100
rect 13132 23154 13524 23156
rect 13132 23102 13246 23154
rect 13298 23102 13524 23154
rect 13132 23100 13524 23102
rect 10332 23044 10388 23054
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 10332 22596 10388 22988
rect 10332 22530 10388 22540
rect 12460 23042 12516 23054
rect 12460 22990 12462 23042
rect 12514 22990 12516 23042
rect 12460 22594 12516 22990
rect 12460 22542 12462 22594
rect 12514 22542 12516 22594
rect 12460 22530 12516 22542
rect 12572 22820 12628 22830
rect 12572 22260 12628 22764
rect 12572 22258 12740 22260
rect 12572 22206 12574 22258
rect 12626 22206 12740 22258
rect 12572 22204 12740 22206
rect 12572 22194 12628 22204
rect 4284 21588 4340 21598
rect 12684 21588 12740 22204
rect 12796 22258 12852 22270
rect 12796 22206 12798 22258
rect 12850 22206 12852 22258
rect 12796 21812 12852 22206
rect 12796 21746 12852 21756
rect 12684 21532 12964 21588
rect 4284 21494 4340 21532
rect 10220 21476 10276 21486
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 10220 20804 10276 21420
rect 12348 21476 12404 21486
rect 12348 21474 12628 21476
rect 12348 21422 12350 21474
rect 12402 21422 12628 21474
rect 12348 21420 12628 21422
rect 12348 21410 12404 21420
rect 12572 21026 12628 21420
rect 12572 20974 12574 21026
rect 12626 20974 12628 21026
rect 12572 20962 12628 20974
rect 12908 21026 12964 21532
rect 13132 21586 13188 23100
rect 13244 23090 13300 23100
rect 13468 22932 13524 23100
rect 13468 22866 13524 22876
rect 13580 23154 13972 23156
rect 13580 23102 13918 23154
rect 13970 23102 13972 23154
rect 13580 23100 13972 23102
rect 13468 22596 13524 22606
rect 13468 21698 13524 22540
rect 13468 21646 13470 21698
rect 13522 21646 13524 21698
rect 13468 21634 13524 21646
rect 13580 22258 13636 23100
rect 13916 23090 13972 23100
rect 13580 22206 13582 22258
rect 13634 22206 13636 22258
rect 13132 21534 13134 21586
rect 13186 21534 13188 21586
rect 13132 21522 13188 21534
rect 12908 20974 12910 21026
rect 12962 20974 12964 21026
rect 12908 20962 12964 20974
rect 13580 20916 13636 22206
rect 13580 20850 13636 20860
rect 13692 22146 13748 22158
rect 13692 22094 13694 22146
rect 13746 22094 13748 22146
rect 13692 21810 13748 22094
rect 13692 21758 13694 21810
rect 13746 21758 13748 21810
rect 10220 20738 10276 20748
rect 13468 20804 13524 20814
rect 13468 20710 13524 20748
rect 13692 20802 13748 21758
rect 13804 21812 13860 21822
rect 13804 21718 13860 21756
rect 14028 21810 14084 23548
rect 14140 23538 14196 23548
rect 14252 23378 14308 24558
rect 14476 23938 14532 24668
rect 15036 24722 15092 24892
rect 15372 24946 15428 25452
rect 15372 24894 15374 24946
rect 15426 24894 15428 24946
rect 15372 24882 15428 24894
rect 16156 25506 16324 25508
rect 16156 25454 16270 25506
rect 16322 25454 16324 25506
rect 16156 25452 16324 25454
rect 16156 24948 16212 25452
rect 16268 25442 16324 25452
rect 17388 25564 17500 25620
rect 16940 25396 16996 25406
rect 16940 25302 16996 25340
rect 16156 24854 16212 24892
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24658 15092 24670
rect 15596 24724 15652 24734
rect 15596 24630 15652 24668
rect 14476 23886 14478 23938
rect 14530 23886 14532 23938
rect 14476 23874 14532 23886
rect 14812 23828 14868 23838
rect 14812 23826 14980 23828
rect 14812 23774 14814 23826
rect 14866 23774 14980 23826
rect 14812 23772 14980 23774
rect 14812 23762 14868 23772
rect 14252 23326 14254 23378
rect 14306 23326 14308 23378
rect 14252 23314 14308 23326
rect 14700 23714 14756 23726
rect 14700 23662 14702 23714
rect 14754 23662 14756 23714
rect 14252 23154 14308 23166
rect 14252 23102 14254 23154
rect 14306 23102 14308 23154
rect 14140 22932 14196 22942
rect 14140 22372 14196 22876
rect 14252 22484 14308 23102
rect 14700 23154 14756 23662
rect 14700 23102 14702 23154
rect 14754 23102 14756 23154
rect 14700 23090 14756 23102
rect 14476 22932 14532 22942
rect 14476 22838 14532 22876
rect 14252 22428 14756 22484
rect 14140 22370 14644 22372
rect 14140 22318 14142 22370
rect 14194 22318 14644 22370
rect 14140 22316 14644 22318
rect 14140 22306 14196 22316
rect 14028 21758 14030 21810
rect 14082 21758 14084 21810
rect 14028 21746 14084 21758
rect 14588 21812 14644 22316
rect 14700 22260 14756 22428
rect 14812 22260 14868 22270
rect 14700 22258 14868 22260
rect 14700 22206 14814 22258
rect 14866 22206 14868 22258
rect 14700 22204 14868 22206
rect 14588 21810 14756 21812
rect 14588 21758 14590 21810
rect 14642 21758 14756 21810
rect 14588 21756 14756 21758
rect 14588 21746 14644 21756
rect 13692 20750 13694 20802
rect 13746 20750 13748 20802
rect 13692 20738 13748 20750
rect 13916 21586 13972 21598
rect 13916 21534 13918 21586
rect 13970 21534 13972 21586
rect 13916 20804 13972 21534
rect 13916 20802 14308 20804
rect 13916 20750 13918 20802
rect 13970 20750 14308 20802
rect 13916 20748 14308 20750
rect 13916 20738 13972 20748
rect 12684 20580 12740 20590
rect 12684 20486 12740 20524
rect 13804 20580 13860 20590
rect 13804 20486 13860 20524
rect 14028 20578 14084 20590
rect 14028 20526 14030 20578
rect 14082 20526 14084 20578
rect 14028 19908 14084 20526
rect 14028 19842 14084 19852
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4172 19282 4228 19292
rect 14252 19348 14308 20748
rect 14700 19572 14756 21756
rect 14812 20132 14868 22204
rect 14924 20916 14980 23772
rect 16940 22482 16996 22494
rect 16940 22430 16942 22482
rect 16994 22430 16996 22482
rect 16604 22148 16660 22158
rect 14924 20850 14980 20860
rect 16380 21700 16436 21710
rect 16044 20804 16100 20814
rect 14812 20066 14868 20076
rect 15596 20132 15652 20142
rect 15260 19908 15316 19918
rect 15148 19852 15260 19908
rect 14700 19516 14868 19572
rect 14700 19348 14756 19358
rect 14252 19346 14756 19348
rect 14252 19294 14254 19346
rect 14306 19294 14702 19346
rect 14754 19294 14756 19346
rect 14252 19292 14756 19294
rect 14252 19282 14308 19292
rect 14700 19282 14756 19292
rect 14028 19236 14084 19246
rect 14028 19234 14196 19236
rect 14028 19182 14030 19234
rect 14082 19182 14196 19234
rect 14028 19180 14196 19182
rect 14028 19170 14084 19180
rect 12908 19122 12964 19134
rect 12908 19070 12910 19122
rect 12962 19070 12964 19122
rect 12572 19012 12628 19022
rect 12236 19010 12628 19012
rect 12236 18958 12574 19010
rect 12626 18958 12628 19010
rect 12236 18956 12628 18958
rect 12236 18562 12292 18956
rect 12572 18946 12628 18956
rect 12908 19012 12964 19070
rect 12908 18946 12964 18956
rect 13692 19012 13748 19022
rect 13692 18918 13748 18956
rect 12236 18510 12238 18562
rect 12290 18510 12292 18562
rect 12236 18498 12292 18510
rect 11564 18452 11620 18462
rect 11564 18358 11620 18396
rect 14028 18452 14084 18462
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17780 1988 17790
rect 1932 17686 1988 17724
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 12460 17668 12516 17678
rect 12460 16770 12516 17612
rect 12460 16718 12462 16770
rect 12514 16718 12516 16770
rect 12460 16706 12516 16718
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 14028 16098 14084 18396
rect 14140 17556 14196 19180
rect 14700 19124 14756 19134
rect 14700 19030 14756 19068
rect 14812 18452 14868 19516
rect 14812 18358 14868 18396
rect 14924 19122 14980 19134
rect 14924 19070 14926 19122
rect 14978 19070 14980 19122
rect 14364 18340 14420 18350
rect 14364 18246 14420 18284
rect 14924 18228 14980 19070
rect 14924 18162 14980 18172
rect 15148 17666 15204 19852
rect 15260 19842 15316 19852
rect 15596 19684 15652 20076
rect 15596 19618 15652 19628
rect 15820 20018 15876 20030
rect 15820 19966 15822 20018
rect 15874 19966 15876 20018
rect 15820 19796 15876 19966
rect 15148 17614 15150 17666
rect 15202 17614 15204 17666
rect 15148 17602 15204 17614
rect 15484 19122 15540 19134
rect 15484 19070 15486 19122
rect 15538 19070 15540 19122
rect 15484 18452 15540 19070
rect 15820 19124 15876 19740
rect 15820 19058 15876 19068
rect 14252 17556 14308 17566
rect 14140 17500 14252 17556
rect 14252 17490 14308 17500
rect 15372 17556 15428 17566
rect 15372 17462 15428 17500
rect 14588 17444 14644 17454
rect 14588 16994 14644 17388
rect 14588 16942 14590 16994
rect 14642 16942 14644 16994
rect 14588 16930 14644 16942
rect 14700 16996 14756 17006
rect 14700 16210 14756 16940
rect 15372 16884 15428 16894
rect 15484 16884 15540 18396
rect 16044 18450 16100 20748
rect 16380 20802 16436 21644
rect 16380 20750 16382 20802
rect 16434 20750 16436 20802
rect 16380 20738 16436 20750
rect 16604 20690 16660 22092
rect 16940 21700 16996 22430
rect 17388 22482 17444 25564
rect 17500 25554 17556 25564
rect 19068 25618 19124 25630
rect 19068 25566 19070 25618
rect 19122 25566 19124 25618
rect 18060 25396 18116 25406
rect 18116 25340 18340 25396
rect 18060 25330 18116 25340
rect 18284 24946 18340 25340
rect 18284 24894 18286 24946
rect 18338 24894 18340 24946
rect 18284 24882 18340 24894
rect 18620 24948 18676 24958
rect 18620 24854 18676 24892
rect 18172 24836 18228 24846
rect 18172 24724 18228 24780
rect 18060 24722 18228 24724
rect 18060 24670 18174 24722
rect 18226 24670 18228 24722
rect 18060 24668 18228 24670
rect 17948 22932 18004 22942
rect 17948 22594 18004 22876
rect 17948 22542 17950 22594
rect 18002 22542 18004 22594
rect 17948 22530 18004 22542
rect 17388 22430 17390 22482
rect 17442 22430 17444 22482
rect 17388 22418 17444 22430
rect 17836 22258 17892 22270
rect 17836 22206 17838 22258
rect 17890 22206 17892 22258
rect 16940 21634 16996 21644
rect 17500 21700 17556 21710
rect 17500 21586 17556 21644
rect 17500 21534 17502 21586
rect 17554 21534 17556 21586
rect 17500 21522 17556 21534
rect 17164 21364 17220 21374
rect 17724 21364 17780 21374
rect 17052 20804 17108 20814
rect 17052 20710 17108 20748
rect 16604 20638 16606 20690
rect 16658 20638 16660 20690
rect 16604 20130 16660 20638
rect 17164 20188 17220 21308
rect 17612 21362 17780 21364
rect 17612 21310 17726 21362
rect 17778 21310 17780 21362
rect 17612 21308 17780 21310
rect 17276 20692 17332 20702
rect 17612 20692 17668 21308
rect 17724 21298 17780 21308
rect 17836 20914 17892 22206
rect 17948 22260 18004 22270
rect 17948 22166 18004 22204
rect 18060 21364 18116 24668
rect 18172 24658 18228 24668
rect 18396 24722 18452 24734
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 18396 23492 18452 24670
rect 19068 24164 19124 25566
rect 19516 25618 19572 26124
rect 19516 25566 19518 25618
rect 19570 25566 19572 25618
rect 19516 25554 19572 25566
rect 20076 25506 20132 26348
rect 20076 25454 20078 25506
rect 20130 25454 20132 25506
rect 20076 25442 20132 25454
rect 20300 26178 20356 26190
rect 20300 26126 20302 26178
rect 20354 26126 20356 26178
rect 19404 25282 19460 25294
rect 19404 25230 19406 25282
rect 19458 25230 19460 25282
rect 19404 24836 19460 25230
rect 19404 24770 19460 24780
rect 19628 25282 19684 25294
rect 19628 25230 19630 25282
rect 19682 25230 19684 25282
rect 19404 24610 19460 24622
rect 19404 24558 19406 24610
rect 19458 24558 19460 24610
rect 19180 24164 19236 24174
rect 19068 24162 19236 24164
rect 19068 24110 19182 24162
rect 19234 24110 19236 24162
rect 19068 24108 19236 24110
rect 18956 23828 19012 23838
rect 17836 20862 17838 20914
rect 17890 20862 17892 20914
rect 17836 20850 17892 20862
rect 17948 21362 18116 21364
rect 17948 21310 18062 21362
rect 18114 21310 18116 21362
rect 17948 21308 18116 21310
rect 17276 20690 17612 20692
rect 17276 20638 17278 20690
rect 17330 20638 17612 20690
rect 17276 20636 17612 20638
rect 17276 20626 17332 20636
rect 17612 20598 17668 20636
rect 17836 20578 17892 20590
rect 17836 20526 17838 20578
rect 17890 20526 17892 20578
rect 17164 20132 17444 20188
rect 16604 20078 16606 20130
rect 16658 20078 16660 20130
rect 16604 20066 16660 20078
rect 17388 20130 17444 20132
rect 17388 20078 17390 20130
rect 17442 20078 17444 20130
rect 17388 20066 17444 20078
rect 17724 20130 17780 20142
rect 17724 20078 17726 20130
rect 17778 20078 17780 20130
rect 17724 20020 17780 20078
rect 17724 19954 17780 19964
rect 16492 19796 16548 19806
rect 16492 19702 16548 19740
rect 17724 19348 17780 19358
rect 16044 18398 16046 18450
rect 16098 18398 16100 18450
rect 16044 18340 16100 18398
rect 16044 18274 16100 18284
rect 16268 18562 16324 18574
rect 16268 18510 16270 18562
rect 16322 18510 16324 18562
rect 16268 18228 16324 18510
rect 17724 18450 17780 19292
rect 17836 18676 17892 20526
rect 17948 19236 18004 21308
rect 18060 21298 18116 21308
rect 18284 23436 18900 23492
rect 18172 20804 18228 20814
rect 18284 20804 18340 23436
rect 18844 23378 18900 23436
rect 18844 23326 18846 23378
rect 18898 23326 18900 23378
rect 18844 23314 18900 23326
rect 18396 23268 18452 23278
rect 18396 23174 18452 23212
rect 18508 23156 18564 23166
rect 18956 23156 19012 23772
rect 19068 23268 19124 24108
rect 19180 24098 19236 24108
rect 19404 23826 19460 24558
rect 19404 23774 19406 23826
rect 19458 23774 19460 23826
rect 19292 23716 19348 23726
rect 19292 23622 19348 23660
rect 19068 23202 19124 23212
rect 18508 23062 18564 23100
rect 18732 23100 19012 23156
rect 19180 23156 19236 23166
rect 18508 22258 18564 22270
rect 18508 22206 18510 22258
rect 18562 22206 18564 22258
rect 18396 22146 18452 22158
rect 18396 22094 18398 22146
rect 18450 22094 18452 22146
rect 18396 21812 18452 22094
rect 18396 21364 18452 21756
rect 18396 21298 18452 21308
rect 18508 21586 18564 22206
rect 18508 21534 18510 21586
rect 18562 21534 18564 21586
rect 18172 20802 18340 20804
rect 18172 20750 18174 20802
rect 18226 20750 18340 20802
rect 18172 20748 18340 20750
rect 18172 20738 18228 20748
rect 18172 20244 18228 20282
rect 18172 20178 18228 20188
rect 18172 20020 18228 20030
rect 18060 19908 18116 19918
rect 18060 19814 18116 19852
rect 17948 19170 18004 19180
rect 17948 18676 18004 18686
rect 17836 18674 18004 18676
rect 17836 18622 17950 18674
rect 18002 18622 18004 18674
rect 17836 18620 18004 18622
rect 17948 18564 18004 18620
rect 18172 18674 18228 19964
rect 18172 18622 18174 18674
rect 18226 18622 18228 18674
rect 18172 18610 18228 18622
rect 18060 18564 18116 18574
rect 17948 18508 18060 18564
rect 18060 18498 18116 18508
rect 18284 18564 18340 20748
rect 18508 20804 18564 21534
rect 18620 20916 18676 20926
rect 18620 20822 18676 20860
rect 18508 20738 18564 20748
rect 18732 20188 18788 23100
rect 19180 23062 19236 23100
rect 19404 22148 19460 23774
rect 19628 23828 19684 25230
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20300 25060 20356 26126
rect 20412 25620 20468 25630
rect 20412 25526 20468 25564
rect 20300 25004 20468 25060
rect 20188 24836 20244 24846
rect 20188 24742 20244 24780
rect 20300 24834 20356 24846
rect 20300 24782 20302 24834
rect 20354 24782 20356 24834
rect 19852 24724 19908 24734
rect 19852 24630 19908 24668
rect 20300 24052 20356 24782
rect 20412 24724 20468 25004
rect 20524 24948 20580 24958
rect 20636 24948 20692 26348
rect 20748 26962 20804 26974
rect 20748 26910 20750 26962
rect 20802 26910 20804 26962
rect 20748 25732 20804 26910
rect 21756 26852 21812 27020
rect 22092 26964 22148 26974
rect 22092 26870 22148 26908
rect 23996 26852 24052 26862
rect 21756 26292 21812 26796
rect 23884 26796 23996 26852
rect 21868 26292 21924 26302
rect 21756 26290 21924 26292
rect 21756 26238 21870 26290
rect 21922 26238 21924 26290
rect 21756 26236 21924 26238
rect 21868 26226 21924 26236
rect 22540 26180 22596 26190
rect 22540 26178 22820 26180
rect 22540 26126 22542 26178
rect 22594 26126 22820 26178
rect 22540 26124 22820 26126
rect 22540 26114 22596 26124
rect 20748 25666 20804 25676
rect 22764 25730 22820 26124
rect 22764 25678 22766 25730
rect 22818 25678 22820 25730
rect 22764 25666 22820 25678
rect 23100 25732 23156 25742
rect 23100 25506 23156 25676
rect 23100 25454 23102 25506
rect 23154 25454 23156 25506
rect 23100 25442 23156 25454
rect 23436 25508 23492 25518
rect 22652 25396 22708 25406
rect 20524 24946 20692 24948
rect 20524 24894 20526 24946
rect 20578 24894 20692 24946
rect 20524 24892 20692 24894
rect 22204 25394 22708 25396
rect 22204 25342 22654 25394
rect 22706 25342 22708 25394
rect 22204 25340 22708 25342
rect 22204 24948 22260 25340
rect 22652 25330 22708 25340
rect 23324 25396 23380 25406
rect 23324 25302 23380 25340
rect 22764 25284 22820 25294
rect 22764 25190 22820 25228
rect 20524 24882 20580 24892
rect 20636 24724 20692 24734
rect 20412 24668 20636 24724
rect 20188 23996 20356 24052
rect 20076 23940 20132 23950
rect 20076 23846 20132 23884
rect 19628 23762 19684 23772
rect 20188 23716 20244 23996
rect 20412 23940 20468 23950
rect 20300 23828 20356 23838
rect 20300 23734 20356 23772
rect 19516 23604 19572 23614
rect 19516 23044 19572 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19516 22978 19572 22988
rect 19628 23266 19684 23278
rect 19628 23214 19630 23266
rect 19682 23214 19684 23266
rect 18956 22092 19460 22148
rect 19516 22148 19572 22158
rect 18844 21252 18900 21262
rect 18844 20692 18900 21196
rect 18956 20804 19012 22092
rect 19516 22054 19572 22092
rect 19628 21588 19684 23214
rect 19852 23268 19908 23278
rect 19852 23154 19908 23212
rect 19852 23102 19854 23154
rect 19906 23102 19908 23154
rect 19852 23090 19908 23102
rect 20188 23044 20244 23660
rect 20300 23380 20356 23390
rect 20300 23322 20356 23324
rect 20300 23270 20302 23322
rect 20354 23270 20356 23322
rect 20300 23258 20356 23270
rect 20412 23266 20468 23884
rect 20636 23938 20692 24668
rect 20636 23886 20638 23938
rect 20690 23886 20692 23938
rect 20636 23874 20692 23886
rect 20748 23940 20804 23950
rect 20748 23846 20804 23884
rect 20412 23214 20414 23266
rect 20466 23214 20468 23266
rect 20412 23156 20468 23214
rect 20188 22370 20244 22988
rect 20188 22318 20190 22370
rect 20242 22318 20244 22370
rect 20188 22306 20244 22318
rect 20300 23100 20468 23156
rect 20748 23324 21028 23380
rect 19852 22148 19908 22158
rect 19852 22146 20244 22148
rect 19852 22094 19854 22146
rect 19906 22094 20244 22146
rect 19852 22092 20244 22094
rect 19852 22082 19908 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 22092
rect 20300 22036 20356 23100
rect 20412 22930 20468 22942
rect 20412 22878 20414 22930
rect 20466 22878 20468 22930
rect 20412 22260 20468 22878
rect 20412 22194 20468 22204
rect 20524 22148 20580 22158
rect 20748 22148 20804 23324
rect 20972 23266 21028 23324
rect 20972 23214 20974 23266
rect 21026 23214 21028 23266
rect 20972 23202 21028 23214
rect 20524 22146 20692 22148
rect 20524 22094 20526 22146
rect 20578 22094 20692 22146
rect 20524 22092 20692 22094
rect 20524 22082 20580 22092
rect 20300 21980 20468 22036
rect 19964 21756 20244 21812
rect 19852 21700 19908 21710
rect 19852 21606 19908 21644
rect 18956 20710 19012 20748
rect 19516 20804 19572 20814
rect 19628 20804 19684 21532
rect 19516 20802 19684 20804
rect 19516 20750 19518 20802
rect 19570 20750 19684 20802
rect 19516 20748 19684 20750
rect 18844 20598 18900 20636
rect 18732 20132 18900 20188
rect 18732 20018 18788 20030
rect 18732 19966 18734 20018
rect 18786 19966 18788 20018
rect 18396 19908 18452 19918
rect 18396 19814 18452 19852
rect 18620 19684 18676 19694
rect 18508 19628 18620 19684
rect 18284 18562 18452 18564
rect 18284 18510 18286 18562
rect 18338 18510 18452 18562
rect 18284 18508 18452 18510
rect 18284 18498 18340 18508
rect 17724 18398 17726 18450
rect 17778 18398 17780 18450
rect 17724 18386 17780 18398
rect 16268 18162 16324 18172
rect 16828 18340 16884 18350
rect 15708 17780 15764 17790
rect 16156 17780 16212 17790
rect 15708 17778 16212 17780
rect 15708 17726 15710 17778
rect 15762 17726 16158 17778
rect 16210 17726 16212 17778
rect 15708 17724 16212 17726
rect 15708 17714 15764 17724
rect 16156 17714 16212 17724
rect 15596 17668 15652 17678
rect 15596 17574 15652 17612
rect 16380 17668 16436 17678
rect 15708 17442 15764 17454
rect 15708 17390 15710 17442
rect 15762 17390 15764 17442
rect 15708 17220 15764 17390
rect 16268 17444 16324 17454
rect 16268 17350 16324 17388
rect 16380 17442 16436 17612
rect 16380 17390 16382 17442
rect 16434 17390 16436 17442
rect 15708 17154 15764 17164
rect 15820 16884 15876 16894
rect 15372 16882 15820 16884
rect 15372 16830 15374 16882
rect 15426 16830 15820 16882
rect 15372 16828 15820 16830
rect 15372 16818 15428 16828
rect 15820 16790 15876 16828
rect 16156 16884 16212 16894
rect 16380 16884 16436 17390
rect 16156 16882 16436 16884
rect 16156 16830 16158 16882
rect 16210 16830 16436 16882
rect 16156 16828 16436 16830
rect 16492 17108 16548 17118
rect 16492 16882 16548 17052
rect 16604 16996 16660 17006
rect 16604 16902 16660 16940
rect 16492 16830 16494 16882
rect 16546 16830 16548 16882
rect 14700 16158 14702 16210
rect 14754 16158 14756 16210
rect 14700 16146 14756 16158
rect 14028 16046 14030 16098
rect 14082 16046 14084 16098
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14028 13746 14084 16046
rect 16156 14530 16212 16828
rect 16492 16818 16548 16830
rect 16828 16882 16884 18284
rect 18060 18340 18116 18350
rect 18060 18246 18116 18284
rect 18396 17554 18452 18508
rect 18508 18562 18564 19628
rect 18620 19618 18676 19628
rect 18732 19348 18788 19966
rect 18732 19282 18788 19292
rect 18508 18510 18510 18562
rect 18562 18510 18564 18562
rect 18508 18498 18564 18510
rect 18844 17780 18900 20132
rect 19068 19236 19124 19246
rect 18620 17724 18900 17780
rect 18956 19124 19012 19134
rect 18620 17668 18676 17724
rect 18396 17502 18398 17554
rect 18450 17502 18452 17554
rect 18396 17490 18452 17502
rect 18508 17666 18676 17668
rect 18508 17614 18622 17666
rect 18674 17614 18676 17666
rect 18508 17612 18676 17614
rect 17612 17220 17668 17230
rect 17276 17108 17332 17118
rect 17500 17108 17556 17118
rect 17276 17014 17332 17052
rect 17388 17106 17556 17108
rect 17388 17054 17502 17106
rect 17554 17054 17556 17106
rect 17388 17052 17556 17054
rect 16828 16830 16830 16882
rect 16882 16830 16884 16882
rect 16828 16818 16884 16830
rect 16156 14478 16158 14530
rect 16210 14478 16212 14530
rect 16156 14466 16212 14478
rect 16828 16212 16884 16222
rect 17388 16212 17444 17052
rect 17500 17042 17556 17052
rect 17612 16994 17668 17164
rect 17612 16942 17614 16994
rect 17666 16942 17668 16994
rect 17612 16930 17668 16942
rect 16828 16210 17444 16212
rect 16828 16158 16830 16210
rect 16882 16158 17444 16210
rect 16828 16156 17444 16158
rect 17500 16884 17556 16894
rect 17500 16212 17556 16828
rect 18508 16772 18564 17612
rect 18620 17602 18676 17612
rect 18844 17556 18900 17566
rect 18956 17556 19012 19068
rect 19068 18450 19124 19180
rect 19516 18788 19572 20748
rect 19852 20580 19908 20590
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 18386 19124 18398
rect 19292 18732 19572 18788
rect 19628 20578 19908 20580
rect 19628 20526 19854 20578
rect 19906 20526 19908 20578
rect 19628 20524 19908 20526
rect 19964 20580 20020 21756
rect 20300 21588 20356 21598
rect 20188 21586 20356 21588
rect 20188 21534 20302 21586
rect 20354 21534 20356 21586
rect 20188 21532 20356 21534
rect 20076 20804 20132 20814
rect 20188 20804 20244 21532
rect 20300 21522 20356 21532
rect 20132 20748 20244 20804
rect 20412 21476 20468 21980
rect 20076 20710 20132 20748
rect 19964 20524 20244 20580
rect 19292 18340 19348 18732
rect 19292 18274 19348 18284
rect 19404 18564 19460 18574
rect 19628 18564 19684 20524
rect 19852 20514 19908 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20076 20132 20132 20142
rect 20076 19234 20132 20076
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 20076 19170 20132 19182
rect 20188 19236 20244 20524
rect 20412 20244 20468 21420
rect 20524 21812 20580 21822
rect 20524 20802 20580 21756
rect 20636 21700 20692 22092
rect 20636 21634 20692 21644
rect 20524 20750 20526 20802
rect 20578 20750 20580 20802
rect 20524 20738 20580 20750
rect 20636 20692 20692 20702
rect 20748 20692 20804 22092
rect 20860 23154 20916 23166
rect 20860 23102 20862 23154
rect 20914 23102 20916 23154
rect 20860 21252 20916 23102
rect 21308 23156 21364 23166
rect 20972 22930 21028 22942
rect 20972 22878 20974 22930
rect 21026 22878 21028 22930
rect 20972 21364 21028 22878
rect 21308 22596 21364 23100
rect 21084 22594 21364 22596
rect 21084 22542 21310 22594
rect 21362 22542 21364 22594
rect 21084 22540 21364 22542
rect 21084 21698 21140 22540
rect 21308 22530 21364 22540
rect 21644 23156 21700 23166
rect 21644 22594 21700 23100
rect 21644 22542 21646 22594
rect 21698 22542 21700 22594
rect 21532 22146 21588 22158
rect 21532 22094 21534 22146
rect 21586 22094 21588 22146
rect 21084 21646 21086 21698
rect 21138 21646 21140 21698
rect 21084 21634 21140 21646
rect 21308 22036 21364 22046
rect 21308 21474 21364 21980
rect 21308 21422 21310 21474
rect 21362 21422 21364 21474
rect 21308 21410 21364 21422
rect 21532 21476 21588 22094
rect 21532 21410 21588 21420
rect 20972 21298 21028 21308
rect 20860 21186 20916 21196
rect 20636 20690 20804 20692
rect 20636 20638 20638 20690
rect 20690 20638 20804 20690
rect 20636 20636 20804 20638
rect 20860 21028 20916 21038
rect 20860 20802 20916 20972
rect 20860 20750 20862 20802
rect 20914 20750 20916 20802
rect 20636 20626 20692 20636
rect 20412 20178 20468 20188
rect 20860 20188 20916 20750
rect 21644 20802 21700 22542
rect 22204 22370 22260 24892
rect 23324 23380 23380 23390
rect 23436 23380 23492 25452
rect 23772 25284 23828 25294
rect 23772 25190 23828 25228
rect 23884 23940 23940 26796
rect 23996 26786 24052 26796
rect 23996 26180 24052 26190
rect 23996 25394 24052 26124
rect 23996 25342 23998 25394
rect 24050 25342 24052 25394
rect 23996 25330 24052 25342
rect 24108 25508 24164 25518
rect 24108 25394 24164 25452
rect 24108 25342 24110 25394
rect 24162 25342 24164 25394
rect 24108 25284 24164 25342
rect 24220 25396 24276 27134
rect 24668 26962 24724 26974
rect 24668 26910 24670 26962
rect 24722 26910 24724 26962
rect 24668 26852 24724 26910
rect 25228 26852 25284 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 39788 36372 39844 36382
rect 39788 36278 39844 36316
rect 40236 36258 40292 36270
rect 40236 36206 40238 36258
rect 40290 36206 40292 36258
rect 40236 35700 40292 36206
rect 40236 35634 40292 35644
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 24668 26786 24724 26796
rect 24780 26796 25284 26852
rect 25340 26852 25396 26862
rect 24668 26180 24724 26190
rect 24780 26180 24836 26796
rect 25340 26514 25396 26796
rect 25340 26462 25342 26514
rect 25394 26462 25396 26514
rect 25340 26450 25396 26462
rect 24724 26124 24836 26180
rect 24668 26086 24724 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 24220 25330 24276 25340
rect 37660 25506 37716 25518
rect 37660 25454 37662 25506
rect 37714 25454 37716 25506
rect 24108 25218 24164 25228
rect 25116 25284 25172 25294
rect 25172 25228 25284 25284
rect 25116 25218 25172 25228
rect 24444 24836 24500 24846
rect 23324 23378 23492 23380
rect 23324 23326 23326 23378
rect 23378 23326 23492 23378
rect 23324 23324 23492 23326
rect 23548 23938 23940 23940
rect 23548 23886 23886 23938
rect 23938 23886 23940 23938
rect 23548 23884 23940 23886
rect 23324 23314 23380 23324
rect 22988 23156 23044 23166
rect 22988 23062 23044 23100
rect 23436 23156 23492 23166
rect 22204 22318 22206 22370
rect 22258 22318 22260 22370
rect 22092 22260 22148 22270
rect 22092 22166 22148 22204
rect 21868 22148 21924 22158
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20738 21700 20750
rect 21756 22146 21924 22148
rect 21756 22094 21870 22146
rect 21922 22094 21924 22146
rect 21756 22092 21924 22094
rect 21756 20188 21812 22092
rect 21868 22082 21924 22092
rect 22204 22036 22260 22318
rect 22764 22260 22820 22270
rect 22764 22166 22820 22204
rect 22204 21970 22260 21980
rect 23100 22146 23156 22158
rect 23100 22094 23102 22146
rect 23154 22094 23156 22146
rect 23100 21812 23156 22094
rect 23100 21746 23156 21756
rect 23436 21810 23492 23100
rect 23548 22372 23604 23884
rect 23884 23874 23940 23884
rect 24332 24834 24500 24836
rect 24332 24782 24446 24834
rect 24498 24782 24500 24834
rect 24332 24780 24500 24782
rect 24332 23156 24388 24780
rect 24444 24770 24500 24780
rect 24556 24724 24612 24734
rect 24556 24630 24612 24668
rect 25228 24722 25284 25228
rect 25228 24670 25230 24722
rect 25282 24670 25284 24722
rect 24444 24500 24500 24510
rect 24444 24498 24724 24500
rect 24444 24446 24446 24498
rect 24498 24446 24724 24498
rect 24444 24444 24724 24446
rect 24444 24434 24500 24444
rect 24668 24050 24724 24444
rect 24668 23998 24670 24050
rect 24722 23998 24724 24050
rect 24668 23986 24724 23998
rect 25228 23266 25284 24670
rect 25340 24834 25396 24846
rect 25340 24782 25342 24834
rect 25394 24782 25396 24834
rect 25340 24052 25396 24782
rect 25564 24724 25620 24734
rect 25564 24630 25620 24668
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 25340 23986 25396 23996
rect 26796 24052 26852 24062
rect 26796 23958 26852 23996
rect 37660 24052 37716 25454
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 37660 23986 37716 23996
rect 27244 23714 27300 23726
rect 27244 23662 27246 23714
rect 27298 23662 27300 23714
rect 25228 23214 25230 23266
rect 25282 23214 25284 23266
rect 25228 23202 25284 23214
rect 25340 23268 25396 23278
rect 25340 23266 25508 23268
rect 25340 23214 25342 23266
rect 25394 23214 25508 23266
rect 25340 23212 25508 23214
rect 25340 23202 25396 23212
rect 24332 23090 24388 23100
rect 23548 22278 23604 22316
rect 24332 22932 24388 22942
rect 24220 22260 24276 22270
rect 23436 21758 23438 21810
rect 23490 21758 23492 21810
rect 23436 21746 23492 21758
rect 23996 22258 24276 22260
rect 23996 22206 24222 22258
rect 24274 22206 24276 22258
rect 23996 22204 24276 22206
rect 23996 21810 24052 22204
rect 24220 22194 24276 22204
rect 23996 21758 23998 21810
rect 24050 21758 24052 21810
rect 23996 21746 24052 21758
rect 24108 21812 24164 21822
rect 21980 21700 22036 21710
rect 20860 20132 21140 20188
rect 20636 19236 20692 19246
rect 20188 19180 20636 19236
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19404 18562 19684 18564
rect 19404 18510 19406 18562
rect 19458 18510 19684 18562
rect 19404 18508 19684 18510
rect 19404 18452 19460 18508
rect 19404 17892 19460 18396
rect 19964 18450 20020 18462
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19404 17826 19460 17836
rect 19516 18338 19572 18350
rect 19516 18286 19518 18338
rect 19570 18286 19572 18338
rect 18844 17554 19012 17556
rect 18844 17502 18846 17554
rect 18898 17502 19012 17554
rect 18844 17500 19012 17502
rect 18844 17490 18900 17500
rect 18732 17442 18788 17454
rect 18732 17390 18734 17442
rect 18786 17390 18788 17442
rect 18732 17220 18788 17390
rect 18732 17154 18788 17164
rect 19516 17108 19572 18286
rect 19964 18340 20020 18398
rect 20636 18450 20692 19180
rect 20636 18398 20638 18450
rect 20690 18398 20692 18450
rect 20636 18386 20692 18398
rect 19964 18274 20020 18284
rect 20972 18340 21028 18350
rect 20972 18246 21028 18284
rect 20524 18226 20580 18238
rect 20524 18174 20526 18226
rect 20578 18174 20580 18226
rect 19852 17668 19908 17678
rect 19908 17612 20020 17668
rect 19852 17574 19908 17612
rect 19852 17444 19908 17454
rect 19516 17042 19572 17052
rect 19628 17442 19908 17444
rect 19628 17390 19854 17442
rect 19906 17390 19908 17442
rect 19628 17388 19908 17390
rect 18508 16706 18564 16716
rect 18620 16884 18676 16894
rect 17500 16210 17892 16212
rect 17500 16158 17502 16210
rect 17554 16158 17892 16210
rect 17500 16156 17892 16158
rect 16492 14418 16548 14430
rect 16492 14366 16494 14418
rect 16546 14366 16548 14418
rect 14700 14308 14756 14318
rect 14700 13858 14756 14252
rect 16380 14308 16436 14318
rect 16380 14214 16436 14252
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13682 14084 13694
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 16492 13188 16548 14366
rect 16828 13860 16884 16156
rect 17500 15538 17556 16156
rect 17500 15486 17502 15538
rect 17554 15486 17556 15538
rect 17500 15474 17556 15486
rect 17836 16098 17892 16156
rect 18620 16210 18676 16828
rect 19628 16884 19684 17388
rect 19852 17378 19908 17388
rect 19964 17444 20020 17612
rect 19964 17378 20020 17388
rect 20188 17666 20244 17678
rect 20188 17614 20190 17666
rect 20242 17614 20244 17666
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 17106 20244 17614
rect 20188 17054 20190 17106
rect 20242 17054 20244 17106
rect 20188 17042 20244 17054
rect 20412 17554 20468 17566
rect 20412 17502 20414 17554
rect 20466 17502 20468 17554
rect 20412 17108 20468 17502
rect 20412 17042 20468 17052
rect 20076 16996 20132 17006
rect 20524 16996 20580 18174
rect 20860 18228 20916 18238
rect 20860 18134 20916 18172
rect 20636 17668 20692 17678
rect 20636 17574 20692 17612
rect 20748 17444 20804 17454
rect 20804 17388 20916 17444
rect 20748 17378 20804 17388
rect 20748 17220 20804 17230
rect 20524 16940 20692 16996
rect 20076 16902 20132 16940
rect 19628 16818 19684 16828
rect 20300 16884 20356 16894
rect 20300 16790 20356 16828
rect 18620 16158 18622 16210
rect 18674 16158 18676 16210
rect 18620 16146 18676 16158
rect 19180 16772 19236 16782
rect 17836 16046 17838 16098
rect 17890 16046 17892 16098
rect 17836 15148 17892 16046
rect 17836 15092 18004 15148
rect 17948 14644 18004 15092
rect 17612 14642 18004 14644
rect 17612 14590 17950 14642
rect 18002 14590 18004 14642
rect 17612 14588 18004 14590
rect 16492 13122 16548 13132
rect 16716 13804 16884 13860
rect 17164 14306 17220 14318
rect 17164 14254 17166 14306
rect 17218 14254 17220 14306
rect 16716 12628 16772 13804
rect 16828 13634 16884 13646
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 16828 13412 16884 13582
rect 17164 13412 17220 14254
rect 17500 14306 17556 14318
rect 17500 14254 17502 14306
rect 17554 14254 17556 14306
rect 17388 13860 17444 13870
rect 16828 13356 17332 13412
rect 17164 13188 17220 13198
rect 17164 13074 17220 13132
rect 17164 13022 17166 13074
rect 17218 13022 17220 13074
rect 17164 13010 17220 13022
rect 17164 12852 17220 12862
rect 17276 12852 17332 13356
rect 17388 13186 17444 13804
rect 17388 13134 17390 13186
rect 17442 13134 17444 13186
rect 17388 13122 17444 13134
rect 17164 12850 17332 12852
rect 17164 12798 17166 12850
rect 17218 12798 17332 12850
rect 17164 12796 17332 12798
rect 17164 12786 17220 12796
rect 16716 12572 17108 12628
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 16828 5236 16884 5246
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16828 800 16884 5180
rect 17052 5122 17108 12572
rect 17052 5070 17054 5122
rect 17106 5070 17108 5122
rect 17052 5058 17108 5070
rect 17276 4450 17332 12796
rect 17276 4398 17278 4450
rect 17330 4398 17332 4450
rect 17276 4386 17332 4398
rect 17500 3556 17556 14254
rect 17612 13746 17668 14588
rect 17612 13694 17614 13746
rect 17666 13694 17668 13746
rect 17612 13682 17668 13694
rect 17948 13074 18004 14588
rect 19180 14530 19236 16716
rect 20524 16772 20580 16782
rect 20524 16678 20580 16716
rect 20076 16660 20132 16670
rect 20076 15876 20132 16604
rect 20076 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20076 15428 20132 15438
rect 20188 15428 20244 15820
rect 20076 15426 20244 15428
rect 20076 15374 20078 15426
rect 20130 15374 20244 15426
rect 20076 15372 20244 15374
rect 20636 15428 20692 16940
rect 20748 16882 20804 17164
rect 20748 16830 20750 16882
rect 20802 16830 20804 16882
rect 20748 16818 20804 16830
rect 20076 15362 20132 15372
rect 20636 15334 20692 15372
rect 20748 16548 20804 16558
rect 20748 16210 20804 16492
rect 20748 16158 20750 16210
rect 20802 16158 20804 16210
rect 20412 15314 20468 15326
rect 20412 15262 20414 15314
rect 20466 15262 20468 15314
rect 19516 15204 19572 15214
rect 19516 14754 19572 15148
rect 20188 15204 20244 15214
rect 20188 15110 20244 15148
rect 19516 14702 19518 14754
rect 19570 14702 19572 14754
rect 19516 14690 19572 14702
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 19180 14466 19236 14478
rect 18284 14308 18340 14318
rect 18284 13858 18340 14252
rect 19404 14308 19460 14318
rect 19404 14214 19460 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 18284 13806 18286 13858
rect 18338 13806 18340 13858
rect 18284 13794 18340 13806
rect 17948 13022 17950 13074
rect 18002 13022 18004 13074
rect 17948 13010 18004 13022
rect 20412 13634 20468 15262
rect 20412 13582 20414 13634
rect 20466 13582 20468 13634
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20412 5906 20468 13582
rect 20412 5854 20414 5906
rect 20466 5854 20468 5906
rect 20412 5842 20468 5854
rect 20188 5684 20244 5694
rect 18060 5236 18116 5246
rect 18060 5142 18116 5180
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 17612 4450 17668 4462
rect 17612 4398 17614 4450
rect 17666 4398 17668 4450
rect 17612 4340 17668 4398
rect 17724 4340 17780 4350
rect 17612 4338 17780 4340
rect 17612 4286 17726 4338
rect 17778 4286 17780 4338
rect 17612 4284 17780 4286
rect 17724 4274 17780 4284
rect 17724 4116 17780 4126
rect 17612 3556 17668 3566
rect 17500 3554 17668 3556
rect 17500 3502 17614 3554
rect 17666 3502 17668 3554
rect 17500 3500 17668 3502
rect 17612 3490 17668 3500
rect 17724 3388 17780 4060
rect 18732 4116 18788 4126
rect 18732 4022 18788 4060
rect 18620 3666 18676 3678
rect 18620 3614 18622 3666
rect 18674 3614 18676 3666
rect 18620 3388 18676 3614
rect 17500 3332 17780 3388
rect 18172 3332 18676 3388
rect 17500 800 17556 3332
rect 18172 800 18228 3332
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 5628
rect 20748 4340 20804 16158
rect 20860 15540 20916 17388
rect 20972 16772 21028 16782
rect 21084 16772 21140 20132
rect 20972 16770 21140 16772
rect 20972 16718 20974 16770
rect 21026 16718 21140 16770
rect 20972 16716 21140 16718
rect 21308 20132 21812 20188
rect 21868 21698 22036 21700
rect 21868 21646 21982 21698
rect 22034 21646 22036 21698
rect 21868 21644 22036 21646
rect 20972 16706 21028 16716
rect 20972 15540 21028 15550
rect 20860 15538 21028 15540
rect 20860 15486 20974 15538
rect 21026 15486 21028 15538
rect 20860 15484 21028 15486
rect 20972 15474 21028 15484
rect 21308 15540 21364 20132
rect 21420 20020 21476 20030
rect 21420 19234 21476 19964
rect 21420 19182 21422 19234
rect 21474 19182 21476 19234
rect 21420 19170 21476 19182
rect 21532 19908 21588 19918
rect 21420 17892 21476 17902
rect 21532 17892 21588 19852
rect 21868 19908 21924 21644
rect 21980 21634 22036 21644
rect 22764 21700 22820 21710
rect 22204 21588 22260 21598
rect 22204 21494 22260 21532
rect 22764 21588 22820 21644
rect 23324 21698 23380 21710
rect 23324 21646 23326 21698
rect 23378 21646 23380 21698
rect 22764 21586 23044 21588
rect 22764 21534 22766 21586
rect 22818 21534 23044 21586
rect 22764 21532 23044 21534
rect 22764 21522 22820 21532
rect 22764 21364 22820 21374
rect 22316 20802 22372 20814
rect 22316 20750 22318 20802
rect 22370 20750 22372 20802
rect 21868 19842 21924 19852
rect 21980 20578 22036 20590
rect 21980 20526 21982 20578
rect 22034 20526 22036 20578
rect 21980 19796 22036 20526
rect 22316 20132 22372 20750
rect 22316 20038 22372 20076
rect 21980 19730 22036 19740
rect 22092 19460 22148 19470
rect 21868 19458 22148 19460
rect 21868 19406 22094 19458
rect 22146 19406 22148 19458
rect 21868 19404 22148 19406
rect 21756 19236 21812 19246
rect 21756 19142 21812 19180
rect 21420 17890 21588 17892
rect 21420 17838 21422 17890
rect 21474 17838 21588 17890
rect 21420 17836 21588 17838
rect 21644 17892 21700 17902
rect 21420 17220 21476 17836
rect 21644 17798 21700 17836
rect 21420 16660 21476 17164
rect 21868 17668 21924 19404
rect 22092 19394 22148 19404
rect 22764 19234 22820 21308
rect 22764 19182 22766 19234
rect 22818 19182 22820 19234
rect 22764 19124 22820 19182
rect 22988 19236 23044 21532
rect 23100 21586 23156 21598
rect 23100 21534 23102 21586
rect 23154 21534 23156 21586
rect 23100 20020 23156 21534
rect 23100 19954 23156 19964
rect 23324 19684 23380 21646
rect 23884 21586 23940 21598
rect 23884 21534 23886 21586
rect 23938 21534 23940 21586
rect 23884 21028 23940 21534
rect 23884 20962 23940 20972
rect 24108 20188 24164 21756
rect 24332 21810 24388 22876
rect 25340 22932 25396 22942
rect 25340 22838 25396 22876
rect 25452 22484 25508 23212
rect 25564 22484 25620 22494
rect 25452 22428 25564 22484
rect 25564 22418 25620 22428
rect 26348 22484 26404 22494
rect 26348 22390 26404 22428
rect 24332 21758 24334 21810
rect 24386 21758 24388 21810
rect 24332 21746 24388 21758
rect 25228 22372 25284 22382
rect 23884 20132 24164 20188
rect 25228 20914 25284 22316
rect 26796 22372 26852 22382
rect 27244 22372 27300 23662
rect 37660 23154 37716 23166
rect 37660 23102 37662 23154
rect 37714 23102 37716 23154
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 37660 22484 37716 23102
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 37660 22418 37716 22428
rect 26852 22316 27300 22372
rect 26796 22278 26852 22316
rect 25788 21812 25844 21822
rect 25788 21718 25844 21756
rect 26796 21698 26852 21710
rect 26796 21646 26798 21698
rect 26850 21646 26852 21698
rect 25564 21586 25620 21598
rect 25564 21534 25566 21586
rect 25618 21534 25620 21586
rect 25564 21364 25620 21534
rect 26236 21588 26292 21598
rect 26572 21588 26628 21598
rect 26236 21586 26628 21588
rect 26236 21534 26238 21586
rect 26290 21534 26574 21586
rect 26626 21534 26628 21586
rect 26236 21532 26628 21534
rect 26236 21522 26292 21532
rect 26572 21522 26628 21532
rect 26796 21588 26852 21646
rect 26796 21522 26852 21532
rect 26908 21586 26964 21598
rect 26908 21534 26910 21586
rect 26962 21534 26964 21586
rect 25564 21298 25620 21308
rect 25676 21474 25732 21486
rect 25676 21422 25678 21474
rect 25730 21422 25732 21474
rect 25228 20862 25230 20914
rect 25282 20862 25284 20914
rect 23324 19618 23380 19628
rect 23436 19796 23492 19806
rect 23100 19236 23156 19246
rect 22988 19234 23156 19236
rect 22988 19182 23102 19234
rect 23154 19182 23156 19234
rect 22988 19180 23156 19182
rect 22764 19058 22820 19068
rect 22988 19010 23044 19022
rect 22988 18958 22990 19010
rect 23042 18958 23044 19010
rect 22092 18228 22148 18238
rect 21868 16996 21924 17612
rect 21980 18172 22092 18228
rect 21980 17666 22036 18172
rect 22092 18162 22148 18172
rect 22092 17890 22148 17902
rect 22092 17838 22094 17890
rect 22146 17838 22148 17890
rect 22092 17780 22148 17838
rect 22092 17724 22372 17780
rect 21980 17614 21982 17666
rect 22034 17614 22036 17666
rect 21980 17602 22036 17614
rect 22316 17668 22372 17724
rect 22428 17668 22484 17678
rect 22764 17668 22820 17678
rect 22316 17666 22484 17668
rect 22316 17614 22430 17666
rect 22482 17614 22484 17666
rect 22316 17612 22484 17614
rect 22428 17602 22484 17612
rect 22540 17666 22820 17668
rect 22540 17614 22766 17666
rect 22818 17614 22820 17666
rect 22540 17612 22820 17614
rect 22204 17556 22260 17566
rect 22204 17462 22260 17500
rect 22540 17220 22596 17612
rect 22764 17602 22820 17612
rect 22988 17666 23044 18958
rect 22988 17614 22990 17666
rect 23042 17614 23044 17666
rect 22988 17602 23044 17614
rect 22316 17164 22596 17220
rect 22764 17442 22820 17454
rect 22764 17390 22766 17442
rect 22818 17390 22820 17442
rect 22092 17108 22148 17118
rect 22092 17014 22148 17052
rect 22316 17106 22372 17164
rect 22316 17054 22318 17106
rect 22370 17054 22372 17106
rect 22316 17042 22372 17054
rect 21980 16996 22036 17006
rect 21868 16994 22036 16996
rect 21868 16942 21982 16994
rect 22034 16942 22036 16994
rect 21868 16940 22036 16942
rect 21980 16930 22036 16940
rect 21420 16594 21476 16604
rect 22428 16884 22484 16894
rect 21308 15538 21476 15540
rect 21308 15486 21310 15538
rect 21362 15486 21476 15538
rect 21308 15484 21476 15486
rect 21308 15474 21364 15484
rect 20860 15204 20916 15214
rect 20860 13746 20916 15148
rect 21420 14754 21476 15484
rect 21532 15428 21588 15438
rect 21588 15372 21700 15428
rect 21532 15362 21588 15372
rect 21420 14702 21422 14754
rect 21474 14702 21476 14754
rect 21420 14690 21476 14702
rect 21644 14754 21700 15372
rect 21644 14702 21646 14754
rect 21698 14702 21700 14754
rect 21644 14690 21700 14702
rect 22316 14644 22372 14654
rect 21868 14642 22372 14644
rect 21868 14590 22318 14642
rect 22370 14590 22372 14642
rect 21868 14588 22372 14590
rect 21868 14530 21924 14588
rect 22316 14578 22372 14588
rect 21868 14478 21870 14530
rect 21922 14478 21924 14530
rect 21868 14466 21924 14478
rect 22204 14420 22260 14430
rect 22428 14420 22484 16828
rect 22764 16212 22820 17390
rect 23100 17108 23156 19180
rect 23436 19234 23492 19740
rect 23436 19182 23438 19234
rect 23490 19182 23492 19234
rect 23436 19170 23492 19182
rect 23884 19234 23940 20132
rect 24108 20020 24164 20030
rect 24108 19458 24164 19964
rect 24108 19406 24110 19458
rect 24162 19406 24164 19458
rect 24108 19394 24164 19406
rect 25228 20020 25284 20862
rect 25676 20188 25732 21422
rect 25676 20132 26404 20188
rect 26348 20130 26404 20132
rect 26348 20078 26350 20130
rect 26402 20078 26404 20130
rect 26348 20066 26404 20078
rect 25564 20020 25620 20030
rect 25228 20018 25620 20020
rect 25228 19966 25566 20018
rect 25618 19966 25620 20018
rect 25228 19964 25620 19966
rect 24444 19348 24500 19358
rect 24444 19254 24500 19292
rect 23884 19182 23886 19234
rect 23938 19182 23940 19234
rect 23884 18452 23940 19182
rect 24556 19236 24612 19246
rect 24556 18564 24612 19180
rect 25228 19234 25284 19964
rect 25564 19954 25620 19964
rect 26908 19796 26964 21534
rect 28476 21588 28532 21598
rect 28476 19906 28532 21532
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21362 40068 21374
rect 40012 21310 40014 21362
rect 40066 21310 40068 21362
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 40012 20916 40068 21310
rect 40012 20850 40068 20860
rect 37660 20018 37716 20030
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 28476 19854 28478 19906
rect 28530 19854 28532 19906
rect 28476 19842 28532 19854
rect 28924 19906 28980 19918
rect 28924 19854 28926 19906
rect 28978 19854 28980 19906
rect 26684 19740 26908 19796
rect 26012 19348 26068 19358
rect 26012 19254 26068 19292
rect 26572 19348 26628 19358
rect 25228 19182 25230 19234
rect 25282 19182 25284 19234
rect 24556 18498 24612 18508
rect 24668 19122 24724 19134
rect 24668 19070 24670 19122
rect 24722 19070 24724 19122
rect 23884 18386 23940 18396
rect 24668 18340 24724 19070
rect 24668 18274 24724 18284
rect 23100 17042 23156 17052
rect 24780 17668 24836 17678
rect 25228 17668 25284 19182
rect 26572 18674 26628 19292
rect 26572 18622 26574 18674
rect 26626 18622 26628 18674
rect 26572 18610 26628 18622
rect 25900 18564 25956 18574
rect 25900 18470 25956 18508
rect 26684 18564 26740 19740
rect 26908 19730 26964 19740
rect 28140 19348 28196 19358
rect 28140 19254 28196 19292
rect 28588 19012 28644 19022
rect 28924 19012 28980 19854
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 19348 37716 19966
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37660 19282 37716 19292
rect 28588 19010 28980 19012
rect 28588 18958 28590 19010
rect 28642 18958 28980 19010
rect 28588 18956 28980 18958
rect 27020 18564 27076 18574
rect 26684 18562 27076 18564
rect 26684 18510 26686 18562
rect 26738 18510 27022 18562
rect 27074 18510 27076 18562
rect 26684 18508 27076 18510
rect 26684 18498 26740 18508
rect 27020 18498 27076 18508
rect 27132 18564 27188 18574
rect 28588 18564 28644 18956
rect 27132 18562 27300 18564
rect 27132 18510 27134 18562
rect 27186 18510 27300 18562
rect 27132 18508 27300 18510
rect 27132 18498 27188 18508
rect 25340 18452 25396 18462
rect 25340 18358 25396 18396
rect 26348 18450 26404 18462
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 25788 18340 25844 18350
rect 25676 18338 25844 18340
rect 25676 18286 25790 18338
rect 25842 18286 25844 18338
rect 25676 18284 25844 18286
rect 25564 18228 25620 18238
rect 25564 18134 25620 18172
rect 25564 17780 25620 17790
rect 25676 17780 25732 18284
rect 25788 18274 25844 18284
rect 26348 18340 26404 18398
rect 26348 18274 26404 18284
rect 26124 18228 26180 18238
rect 26124 18134 26180 18172
rect 27132 18228 27188 18238
rect 27132 18134 27188 18172
rect 25564 17778 25732 17780
rect 25564 17726 25566 17778
rect 25618 17726 25732 17778
rect 25564 17724 25732 17726
rect 27244 17780 27300 18508
rect 28476 18508 28644 18564
rect 27692 17780 27748 17790
rect 27244 17724 27692 17780
rect 25564 17714 25620 17724
rect 27692 17686 27748 17724
rect 24780 17666 25284 17668
rect 24780 17614 24782 17666
rect 24834 17614 25284 17666
rect 24780 17612 25284 17614
rect 24780 16884 24836 17612
rect 22764 16146 22820 16156
rect 23548 16212 23604 16222
rect 23548 16118 23604 16156
rect 22876 16098 22932 16110
rect 22876 16046 22878 16098
rect 22930 16046 22932 16098
rect 22876 15204 22932 16046
rect 22876 15138 22932 15148
rect 24108 15204 24164 15214
rect 22540 14532 22596 14542
rect 22540 14530 23044 14532
rect 22540 14478 22542 14530
rect 22594 14478 23044 14530
rect 22540 14476 23044 14478
rect 22540 14466 22596 14476
rect 22204 14418 22484 14420
rect 22204 14366 22206 14418
rect 22258 14366 22484 14418
rect 22204 14364 22484 14366
rect 21756 14308 21812 14318
rect 21532 14306 21812 14308
rect 21532 14254 21758 14306
rect 21810 14254 21812 14306
rect 21532 14252 21812 14254
rect 21532 13858 21588 14252
rect 21756 14242 21812 14252
rect 21532 13806 21534 13858
rect 21586 13806 21588 13858
rect 21532 13794 21588 13806
rect 22092 13860 22148 13870
rect 22204 13860 22260 14364
rect 22148 13804 22260 13860
rect 22092 13794 22148 13804
rect 20860 13694 20862 13746
rect 20914 13694 20916 13746
rect 20860 13682 20916 13694
rect 22988 12964 23044 14476
rect 24108 13970 24164 15148
rect 24780 15204 24836 16828
rect 25340 17556 25396 17566
rect 25340 16882 25396 17500
rect 28140 17444 28196 17454
rect 28476 17444 28532 18508
rect 37660 18450 37716 18462
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 37660 17780 37716 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37660 17714 37716 17724
rect 28140 17442 28532 17444
rect 28140 17390 28142 17442
rect 28194 17390 28532 17442
rect 28140 17388 28532 17390
rect 25340 16830 25342 16882
rect 25394 16830 25396 16882
rect 25340 15652 25396 16830
rect 25564 16994 25620 17006
rect 25564 16942 25566 16994
rect 25618 16942 25620 16994
rect 25564 16436 25620 16942
rect 25564 16370 25620 16380
rect 26348 16884 26404 16894
rect 26348 16210 26404 16828
rect 28140 16884 28196 17388
rect 28140 16818 28196 16828
rect 35196 16492 35460 16502
rect 26348 16158 26350 16210
rect 26402 16158 26404 16210
rect 26348 16146 26404 16158
rect 28588 16436 28644 16446
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 25788 15874 25844 15886
rect 25788 15822 25790 15874
rect 25842 15822 25844 15874
rect 25788 15652 25844 15822
rect 25340 15596 25844 15652
rect 25340 15314 25396 15596
rect 25340 15262 25342 15314
rect 25394 15262 25396 15314
rect 25340 15148 25396 15262
rect 24780 15138 24836 15148
rect 24108 13918 24110 13970
rect 24162 13918 24164 13970
rect 24108 13906 24164 13918
rect 25228 15092 25396 15148
rect 25564 15426 25620 15438
rect 25564 15374 25566 15426
rect 25618 15374 25620 15426
rect 23660 13634 23716 13646
rect 23660 13582 23662 13634
rect 23714 13582 23716 13634
rect 23660 12964 23716 13582
rect 22988 12962 23716 12964
rect 22988 12910 22990 12962
rect 23042 12910 23716 12962
rect 22988 12908 23716 12910
rect 22988 12898 23044 12908
rect 23212 12738 23268 12750
rect 23212 12686 23214 12738
rect 23266 12686 23268 12738
rect 23212 10164 23268 12686
rect 23212 10098 23268 10108
rect 21420 5684 21476 5694
rect 21420 5590 21476 5628
rect 21084 4340 21140 4350
rect 20748 4338 21140 4340
rect 20748 4286 21086 4338
rect 21138 4286 21140 4338
rect 20748 4284 21140 4286
rect 21084 4274 21140 4284
rect 20860 4116 20916 4126
rect 20860 800 20916 4060
rect 22092 4116 22148 4126
rect 22092 4022 22148 4060
rect 23660 3554 23716 12908
rect 23772 10164 23828 10174
rect 23772 5122 23828 10108
rect 23996 5236 24052 5246
rect 23772 5070 23774 5122
rect 23826 5070 23828 5122
rect 23772 5058 23828 5070
rect 23884 5180 23996 5236
rect 23660 3502 23662 3554
rect 23714 3502 23716 3554
rect 23660 3490 23716 3502
rect 22204 3442 22260 3454
rect 22204 3390 22206 3442
rect 22258 3390 22260 3442
rect 21084 3332 21140 3342
rect 21084 3330 21588 3332
rect 21084 3278 21086 3330
rect 21138 3278 21588 3330
rect 21084 3276 21588 3278
rect 21084 3266 21140 3276
rect 21532 800 21588 3276
rect 22204 800 22260 3390
rect 22876 3444 22932 3454
rect 23884 3388 23940 5180
rect 23996 5170 24052 5180
rect 24780 5236 24836 5246
rect 24780 5142 24836 5180
rect 25228 5012 25284 15092
rect 25004 4956 25284 5012
rect 22876 800 22932 3388
rect 23660 3332 23940 3388
rect 24892 4116 24948 4126
rect 23660 980 23716 3332
rect 23548 924 23716 980
rect 23548 800 23604 924
rect 24892 800 24948 4060
rect 25004 3554 25060 4956
rect 25564 4338 25620 15374
rect 25564 4286 25566 4338
rect 25618 4286 25620 4338
rect 25564 4274 25620 4286
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 25004 3502 25006 3554
rect 25058 3502 25060 3554
rect 25004 3490 25060 3502
rect 25564 3666 25620 3678
rect 25564 3614 25566 3666
rect 25618 3614 25620 3666
rect 25564 3444 25620 3614
rect 25564 3378 25620 3388
rect 25676 3668 25732 3678
rect 25676 1652 25732 3612
rect 28588 3554 28644 16380
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3490 28644 3502
rect 25564 1596 25732 1652
rect 25564 800 25620 1596
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24864 0 24976 800
rect 25536 0 25648 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 22876 38220 22932 38276
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 24892 37436 24948 37492
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 20412 26962 20468 26964
rect 20412 26910 20414 26962
rect 20414 26910 20466 26962
rect 20466 26910 20468 26962
rect 20412 26908 20468 26910
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 4172 26236 4228 26292
rect 1932 24892 1988 24948
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 20860 1988 20916
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 18172 26178 18228 26180
rect 18172 26126 18174 26178
rect 18174 26126 18226 26178
rect 18226 26126 18228 26178
rect 18172 26124 18228 26126
rect 19516 26124 19572 26180
rect 16268 25564 16324 25620
rect 4284 25506 4340 25508
rect 4284 25454 4286 25506
rect 4286 25454 4338 25506
rect 4338 25454 4340 25506
rect 4284 25452 4340 25454
rect 15372 25452 15428 25508
rect 13580 24892 13636 24948
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 12124 24668 12180 24724
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 15036 24892 15092 24948
rect 14476 24668 14532 24724
rect 14140 23548 14196 23604
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 10332 23042 10388 23044
rect 10332 22990 10334 23042
rect 10334 22990 10386 23042
rect 10386 22990 10388 23042
rect 10332 22988 10388 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 10332 22540 10388 22596
rect 12572 22764 12628 22820
rect 4284 21586 4340 21588
rect 4284 21534 4286 21586
rect 4286 21534 4338 21586
rect 4338 21534 4340 21586
rect 4284 21532 4340 21534
rect 12796 21756 12852 21812
rect 10220 21474 10276 21476
rect 10220 21422 10222 21474
rect 10222 21422 10274 21474
rect 10274 21422 10276 21474
rect 10220 21420 10276 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 13468 22876 13524 22932
rect 13468 22540 13524 22596
rect 13580 20860 13636 20916
rect 10220 20748 10276 20804
rect 13468 20802 13524 20804
rect 13468 20750 13470 20802
rect 13470 20750 13522 20802
rect 13522 20750 13524 20802
rect 13468 20748 13524 20750
rect 13804 21810 13860 21812
rect 13804 21758 13806 21810
rect 13806 21758 13858 21810
rect 13858 21758 13860 21810
rect 13804 21756 13860 21758
rect 17500 25564 17556 25620
rect 16940 25394 16996 25396
rect 16940 25342 16942 25394
rect 16942 25342 16994 25394
rect 16994 25342 16996 25394
rect 16940 25340 16996 25342
rect 16156 24946 16212 24948
rect 16156 24894 16158 24946
rect 16158 24894 16210 24946
rect 16210 24894 16212 24946
rect 16156 24892 16212 24894
rect 15596 24722 15652 24724
rect 15596 24670 15598 24722
rect 15598 24670 15650 24722
rect 15650 24670 15652 24722
rect 15596 24668 15652 24670
rect 14140 22876 14196 22932
rect 14476 22930 14532 22932
rect 14476 22878 14478 22930
rect 14478 22878 14530 22930
rect 14530 22878 14532 22930
rect 14476 22876 14532 22878
rect 12684 20578 12740 20580
rect 12684 20526 12686 20578
rect 12686 20526 12738 20578
rect 12738 20526 12740 20578
rect 12684 20524 12740 20526
rect 13804 20578 13860 20580
rect 13804 20526 13806 20578
rect 13806 20526 13858 20578
rect 13858 20526 13860 20578
rect 13804 20524 13860 20526
rect 14028 19852 14084 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4172 19292 4228 19348
rect 16604 22092 16660 22148
rect 14924 20860 14980 20916
rect 16380 21644 16436 21700
rect 16044 20748 16100 20804
rect 14812 20076 14868 20132
rect 15596 20130 15652 20132
rect 15596 20078 15598 20130
rect 15598 20078 15650 20130
rect 15650 20078 15652 20130
rect 15596 20076 15652 20078
rect 15260 19852 15316 19908
rect 12908 18956 12964 19012
rect 13692 19010 13748 19012
rect 13692 18958 13694 19010
rect 13694 18958 13746 19010
rect 13746 18958 13748 19010
rect 13692 18956 13748 18958
rect 11564 18450 11620 18452
rect 11564 18398 11566 18450
rect 11566 18398 11618 18450
rect 11618 18398 11620 18450
rect 11564 18396 11620 18398
rect 14028 18396 14084 18452
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 12460 17612 12516 17668
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 14700 19122 14756 19124
rect 14700 19070 14702 19122
rect 14702 19070 14754 19122
rect 14754 19070 14756 19122
rect 14700 19068 14756 19070
rect 14812 18450 14868 18452
rect 14812 18398 14814 18450
rect 14814 18398 14866 18450
rect 14866 18398 14868 18450
rect 14812 18396 14868 18398
rect 14364 18338 14420 18340
rect 14364 18286 14366 18338
rect 14366 18286 14418 18338
rect 14418 18286 14420 18338
rect 14364 18284 14420 18286
rect 14924 18172 14980 18228
rect 15596 19628 15652 19684
rect 15820 19740 15876 19796
rect 15820 19068 15876 19124
rect 15484 18396 15540 18452
rect 14252 17500 14308 17556
rect 15372 17554 15428 17556
rect 15372 17502 15374 17554
rect 15374 17502 15426 17554
rect 15426 17502 15428 17554
rect 15372 17500 15428 17502
rect 14588 17388 14644 17444
rect 14700 16940 14756 16996
rect 18060 25340 18116 25396
rect 18620 24946 18676 24948
rect 18620 24894 18622 24946
rect 18622 24894 18674 24946
rect 18674 24894 18676 24946
rect 18620 24892 18676 24894
rect 18172 24780 18228 24836
rect 17948 22876 18004 22932
rect 16940 21644 16996 21700
rect 17500 21644 17556 21700
rect 17164 21308 17220 21364
rect 17052 20802 17108 20804
rect 17052 20750 17054 20802
rect 17054 20750 17106 20802
rect 17106 20750 17108 20802
rect 17052 20748 17108 20750
rect 17948 22258 18004 22260
rect 17948 22206 17950 22258
rect 17950 22206 18002 22258
rect 18002 22206 18004 22258
rect 17948 22204 18004 22206
rect 19404 24780 19460 24836
rect 18956 23772 19012 23828
rect 17612 20690 17668 20692
rect 17612 20638 17614 20690
rect 17614 20638 17666 20690
rect 17666 20638 17668 20690
rect 17612 20636 17668 20638
rect 17724 19964 17780 20020
rect 16492 19794 16548 19796
rect 16492 19742 16494 19794
rect 16494 19742 16546 19794
rect 16546 19742 16548 19794
rect 16492 19740 16548 19742
rect 17724 19292 17780 19348
rect 16044 18284 16100 18340
rect 18396 23266 18452 23268
rect 18396 23214 18398 23266
rect 18398 23214 18450 23266
rect 18450 23214 18452 23266
rect 18396 23212 18452 23214
rect 19292 23714 19348 23716
rect 19292 23662 19294 23714
rect 19294 23662 19346 23714
rect 19346 23662 19348 23714
rect 19292 23660 19348 23662
rect 19068 23212 19124 23268
rect 18508 23154 18564 23156
rect 18508 23102 18510 23154
rect 18510 23102 18562 23154
rect 18562 23102 18564 23154
rect 18508 23100 18564 23102
rect 19180 23154 19236 23156
rect 19180 23102 19182 23154
rect 19182 23102 19234 23154
rect 19234 23102 19236 23154
rect 19180 23100 19236 23102
rect 18396 21756 18452 21812
rect 18396 21308 18452 21364
rect 18172 20242 18228 20244
rect 18172 20190 18174 20242
rect 18174 20190 18226 20242
rect 18226 20190 18228 20242
rect 18172 20188 18228 20190
rect 18172 19964 18228 20020
rect 18060 19906 18116 19908
rect 18060 19854 18062 19906
rect 18062 19854 18114 19906
rect 18114 19854 18116 19906
rect 18060 19852 18116 19854
rect 17948 19180 18004 19236
rect 18060 18508 18116 18564
rect 18620 20914 18676 20916
rect 18620 20862 18622 20914
rect 18622 20862 18674 20914
rect 18674 20862 18676 20914
rect 18620 20860 18676 20862
rect 18508 20748 18564 20804
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20412 25618 20468 25620
rect 20412 25566 20414 25618
rect 20414 25566 20466 25618
rect 20466 25566 20468 25618
rect 20412 25564 20468 25566
rect 20188 24834 20244 24836
rect 20188 24782 20190 24834
rect 20190 24782 20242 24834
rect 20242 24782 20244 24834
rect 20188 24780 20244 24782
rect 19852 24722 19908 24724
rect 19852 24670 19854 24722
rect 19854 24670 19906 24722
rect 19906 24670 19908 24722
rect 19852 24668 19908 24670
rect 22092 26962 22148 26964
rect 22092 26910 22094 26962
rect 22094 26910 22146 26962
rect 22146 26910 22148 26962
rect 22092 26908 22148 26910
rect 21756 26796 21812 26852
rect 23996 26796 24052 26852
rect 20748 25676 20804 25732
rect 23100 25676 23156 25732
rect 23436 25506 23492 25508
rect 23436 25454 23438 25506
rect 23438 25454 23490 25506
rect 23490 25454 23492 25506
rect 23436 25452 23492 25454
rect 23324 25394 23380 25396
rect 23324 25342 23326 25394
rect 23326 25342 23378 25394
rect 23378 25342 23380 25394
rect 23324 25340 23380 25342
rect 22764 25282 22820 25284
rect 22764 25230 22766 25282
rect 22766 25230 22818 25282
rect 22818 25230 22820 25282
rect 22764 25228 22820 25230
rect 22204 24892 22260 24948
rect 20636 24668 20692 24724
rect 20076 23938 20132 23940
rect 20076 23886 20078 23938
rect 20078 23886 20130 23938
rect 20130 23886 20132 23938
rect 20076 23884 20132 23886
rect 19628 23772 19684 23828
rect 20412 23884 20468 23940
rect 20300 23826 20356 23828
rect 20300 23774 20302 23826
rect 20302 23774 20354 23826
rect 20354 23774 20356 23826
rect 20300 23772 20356 23774
rect 20188 23660 20244 23716
rect 19516 23548 19572 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19516 22988 19572 23044
rect 19516 22146 19572 22148
rect 19516 22094 19518 22146
rect 19518 22094 19570 22146
rect 19570 22094 19572 22146
rect 19516 22092 19572 22094
rect 18844 21196 18900 21252
rect 19852 23212 19908 23268
rect 20300 23324 20356 23380
rect 20748 23938 20804 23940
rect 20748 23886 20750 23938
rect 20750 23886 20802 23938
rect 20802 23886 20804 23938
rect 20748 23884 20804 23886
rect 20188 22988 20244 23044
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20412 22204 20468 22260
rect 19852 21698 19908 21700
rect 19852 21646 19854 21698
rect 19854 21646 19906 21698
rect 19906 21646 19908 21698
rect 19852 21644 19908 21646
rect 19628 21532 19684 21588
rect 18956 20802 19012 20804
rect 18956 20750 18958 20802
rect 18958 20750 19010 20802
rect 19010 20750 19012 20802
rect 18956 20748 19012 20750
rect 18844 20690 18900 20692
rect 18844 20638 18846 20690
rect 18846 20638 18898 20690
rect 18898 20638 18900 20690
rect 18844 20636 18900 20638
rect 18396 19906 18452 19908
rect 18396 19854 18398 19906
rect 18398 19854 18450 19906
rect 18450 19854 18452 19906
rect 18396 19852 18452 19854
rect 18620 19628 18676 19684
rect 16268 18172 16324 18228
rect 16828 18284 16884 18340
rect 15596 17666 15652 17668
rect 15596 17614 15598 17666
rect 15598 17614 15650 17666
rect 15650 17614 15652 17666
rect 15596 17612 15652 17614
rect 16380 17612 16436 17668
rect 16268 17442 16324 17444
rect 16268 17390 16270 17442
rect 16270 17390 16322 17442
rect 16322 17390 16324 17442
rect 16268 17388 16324 17390
rect 15708 17164 15764 17220
rect 15820 16882 15876 16884
rect 15820 16830 15822 16882
rect 15822 16830 15874 16882
rect 15874 16830 15876 16882
rect 15820 16828 15876 16830
rect 16492 17052 16548 17108
rect 16604 16994 16660 16996
rect 16604 16942 16606 16994
rect 16606 16942 16658 16994
rect 16658 16942 16660 16994
rect 16604 16940 16660 16942
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 18060 18338 18116 18340
rect 18060 18286 18062 18338
rect 18062 18286 18114 18338
rect 18114 18286 18116 18338
rect 18060 18284 18116 18286
rect 18732 19292 18788 19348
rect 19068 19180 19124 19236
rect 18956 19068 19012 19124
rect 17612 17164 17668 17220
rect 17276 17106 17332 17108
rect 17276 17054 17278 17106
rect 17278 17054 17330 17106
rect 17330 17054 17332 17106
rect 17276 17052 17332 17054
rect 17500 16828 17556 16884
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 20412 21420 20468 21476
rect 19292 18284 19348 18340
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20076 20076 20132 20132
rect 20524 21756 20580 21812
rect 20636 21644 20692 21700
rect 20748 22092 20804 22148
rect 21308 23100 21364 23156
rect 21644 23100 21700 23156
rect 21308 21980 21364 22036
rect 21532 21420 21588 21476
rect 20972 21308 21028 21364
rect 20860 21196 20916 21252
rect 20860 20972 20916 21028
rect 20412 20188 20468 20244
rect 23772 25282 23828 25284
rect 23772 25230 23774 25282
rect 23774 25230 23826 25282
rect 23826 25230 23828 25282
rect 23772 25228 23828 25230
rect 23996 26124 24052 26180
rect 24108 25452 24164 25508
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 39788 36370 39844 36372
rect 39788 36318 39790 36370
rect 39790 36318 39842 36370
rect 39842 36318 39844 36370
rect 39788 36316 39844 36318
rect 40236 35644 40292 35700
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 24668 26796 24724 26852
rect 25340 26796 25396 26852
rect 24668 26178 24724 26180
rect 24668 26126 24670 26178
rect 24670 26126 24722 26178
rect 24722 26126 24724 26178
rect 24668 26124 24724 26126
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 24220 25340 24276 25396
rect 24108 25228 24164 25284
rect 25116 25228 25172 25284
rect 22988 23154 23044 23156
rect 22988 23102 22990 23154
rect 22990 23102 23042 23154
rect 23042 23102 23044 23154
rect 22988 23100 23044 23102
rect 23436 23100 23492 23156
rect 22092 22258 22148 22260
rect 22092 22206 22094 22258
rect 22094 22206 22146 22258
rect 22146 22206 22148 22258
rect 22092 22204 22148 22206
rect 22764 22258 22820 22260
rect 22764 22206 22766 22258
rect 22766 22206 22818 22258
rect 22818 22206 22820 22258
rect 22764 22204 22820 22206
rect 22204 21980 22260 22036
rect 23100 21756 23156 21812
rect 24556 24722 24612 24724
rect 24556 24670 24558 24722
rect 24558 24670 24610 24722
rect 24610 24670 24612 24722
rect 24556 24668 24612 24670
rect 25564 24722 25620 24724
rect 25564 24670 25566 24722
rect 25566 24670 25618 24722
rect 25618 24670 25620 24722
rect 25564 24668 25620 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 25340 23996 25396 24052
rect 26796 24050 26852 24052
rect 26796 23998 26798 24050
rect 26798 23998 26850 24050
rect 26850 23998 26852 24050
rect 26796 23996 26852 23998
rect 40012 24892 40068 24948
rect 37660 23996 37716 24052
rect 24332 23100 24388 23156
rect 23548 22370 23604 22372
rect 23548 22318 23550 22370
rect 23550 22318 23602 22370
rect 23602 22318 23604 22370
rect 23548 22316 23604 22318
rect 24332 22876 24388 22932
rect 24108 21810 24164 21812
rect 24108 21758 24110 21810
rect 24110 21758 24162 21810
rect 24162 21758 24164 21810
rect 24108 21756 24164 21758
rect 20636 19180 20692 19236
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19404 18396 19460 18452
rect 19404 17836 19460 17892
rect 18732 17164 18788 17220
rect 19964 18284 20020 18340
rect 20972 18338 21028 18340
rect 20972 18286 20974 18338
rect 20974 18286 21026 18338
rect 21026 18286 21028 18338
rect 20972 18284 21028 18286
rect 19852 17666 19908 17668
rect 19852 17614 19854 17666
rect 19854 17614 19906 17666
rect 19906 17614 19908 17666
rect 19852 17612 19908 17614
rect 19516 17052 19572 17108
rect 18508 16716 18564 16772
rect 18620 16828 18676 16884
rect 14700 14252 14756 14308
rect 16380 14306 16436 14308
rect 16380 14254 16382 14306
rect 16382 14254 16434 14306
rect 16434 14254 16436 14306
rect 16380 14252 16436 14254
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 19964 17388 20020 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20412 17052 20468 17108
rect 20076 16994 20132 16996
rect 20076 16942 20078 16994
rect 20078 16942 20130 16994
rect 20130 16942 20132 16994
rect 20076 16940 20132 16942
rect 20860 18226 20916 18228
rect 20860 18174 20862 18226
rect 20862 18174 20914 18226
rect 20914 18174 20916 18226
rect 20860 18172 20916 18174
rect 20636 17666 20692 17668
rect 20636 17614 20638 17666
rect 20638 17614 20690 17666
rect 20690 17614 20692 17666
rect 20636 17612 20692 17614
rect 20748 17388 20804 17444
rect 20748 17164 20804 17220
rect 19628 16828 19684 16884
rect 20300 16882 20356 16884
rect 20300 16830 20302 16882
rect 20302 16830 20354 16882
rect 20354 16830 20356 16882
rect 20300 16828 20356 16830
rect 19180 16716 19236 16772
rect 16492 13132 16548 13188
rect 17388 13804 17444 13860
rect 17164 13132 17220 13188
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 16828 5180 16884 5236
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 20524 16770 20580 16772
rect 20524 16718 20526 16770
rect 20526 16718 20578 16770
rect 20578 16718 20580 16770
rect 20524 16716 20580 16718
rect 20076 16604 20132 16660
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20636 15426 20692 15428
rect 20636 15374 20638 15426
rect 20638 15374 20690 15426
rect 20690 15374 20692 15426
rect 20636 15372 20692 15374
rect 20748 16492 20804 16548
rect 19516 15148 19572 15204
rect 20188 15202 20244 15204
rect 20188 15150 20190 15202
rect 20190 15150 20242 15202
rect 20242 15150 20244 15202
rect 20188 15148 20244 15150
rect 18284 14252 18340 14308
rect 19404 14306 19460 14308
rect 19404 14254 19406 14306
rect 19406 14254 19458 14306
rect 19458 14254 19460 14306
rect 19404 14252 19460 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20188 5628 20244 5684
rect 18060 5234 18116 5236
rect 18060 5182 18062 5234
rect 18062 5182 18114 5234
rect 18114 5182 18116 5234
rect 18060 5180 18116 5182
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 17724 4060 17780 4116
rect 18732 4114 18788 4116
rect 18732 4062 18734 4114
rect 18734 4062 18786 4114
rect 18786 4062 18788 4114
rect 18732 4060 18788 4062
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21420 19964 21476 20020
rect 21532 19852 21588 19908
rect 22764 21644 22820 21700
rect 22204 21586 22260 21588
rect 22204 21534 22206 21586
rect 22206 21534 22258 21586
rect 22258 21534 22260 21586
rect 22204 21532 22260 21534
rect 22764 21308 22820 21364
rect 21868 19852 21924 19908
rect 22316 20130 22372 20132
rect 22316 20078 22318 20130
rect 22318 20078 22370 20130
rect 22370 20078 22372 20130
rect 22316 20076 22372 20078
rect 21980 19740 22036 19796
rect 21756 19234 21812 19236
rect 21756 19182 21758 19234
rect 21758 19182 21810 19234
rect 21810 19182 21812 19234
rect 21756 19180 21812 19182
rect 21644 17890 21700 17892
rect 21644 17838 21646 17890
rect 21646 17838 21698 17890
rect 21698 17838 21700 17890
rect 21644 17836 21700 17838
rect 21420 17164 21476 17220
rect 23100 19964 23156 20020
rect 23884 20972 23940 21028
rect 25340 22930 25396 22932
rect 25340 22878 25342 22930
rect 25342 22878 25394 22930
rect 25394 22878 25396 22930
rect 25340 22876 25396 22878
rect 25564 22428 25620 22484
rect 26348 22482 26404 22484
rect 26348 22430 26350 22482
rect 26350 22430 26402 22482
rect 26402 22430 26404 22482
rect 26348 22428 26404 22430
rect 25228 22316 25284 22372
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 37660 22428 37716 22484
rect 26796 22370 26852 22372
rect 26796 22318 26798 22370
rect 26798 22318 26850 22370
rect 26850 22318 26852 22370
rect 26796 22316 26852 22318
rect 25788 21810 25844 21812
rect 25788 21758 25790 21810
rect 25790 21758 25842 21810
rect 25842 21758 25844 21810
rect 25788 21756 25844 21758
rect 26796 21532 26852 21588
rect 25564 21308 25620 21364
rect 23324 19628 23380 19684
rect 23436 19740 23492 19796
rect 22764 19068 22820 19124
rect 21868 17612 21924 17668
rect 22092 18172 22148 18228
rect 22204 17554 22260 17556
rect 22204 17502 22206 17554
rect 22206 17502 22258 17554
rect 22258 17502 22260 17554
rect 22204 17500 22260 17502
rect 22092 17106 22148 17108
rect 22092 17054 22094 17106
rect 22094 17054 22146 17106
rect 22146 17054 22148 17106
rect 22092 17052 22148 17054
rect 21420 16604 21476 16660
rect 22428 16828 22484 16884
rect 20860 15148 20916 15204
rect 21532 15372 21588 15428
rect 24108 19964 24164 20020
rect 24444 19346 24500 19348
rect 24444 19294 24446 19346
rect 24446 19294 24498 19346
rect 24498 19294 24500 19346
rect 24444 19292 24500 19294
rect 24556 19234 24612 19236
rect 24556 19182 24558 19234
rect 24558 19182 24610 19234
rect 24610 19182 24612 19234
rect 24556 19180 24612 19182
rect 28476 21532 28532 21588
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 40012 20860 40068 20916
rect 26908 19740 26964 19796
rect 26012 19346 26068 19348
rect 26012 19294 26014 19346
rect 26014 19294 26066 19346
rect 26066 19294 26068 19346
rect 26012 19292 26068 19294
rect 26572 19292 26628 19348
rect 24556 18508 24612 18564
rect 23884 18396 23940 18452
rect 24668 18284 24724 18340
rect 23100 17052 23156 17108
rect 25900 18562 25956 18564
rect 25900 18510 25902 18562
rect 25902 18510 25954 18562
rect 25954 18510 25956 18562
rect 25900 18508 25956 18510
rect 28140 19346 28196 19348
rect 28140 19294 28142 19346
rect 28142 19294 28194 19346
rect 28194 19294 28196 19346
rect 28140 19292 28196 19294
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 37660 19292 37716 19348
rect 25340 18450 25396 18452
rect 25340 18398 25342 18450
rect 25342 18398 25394 18450
rect 25394 18398 25396 18450
rect 25340 18396 25396 18398
rect 25564 18226 25620 18228
rect 25564 18174 25566 18226
rect 25566 18174 25618 18226
rect 25618 18174 25620 18226
rect 25564 18172 25620 18174
rect 26348 18284 26404 18340
rect 26124 18226 26180 18228
rect 26124 18174 26126 18226
rect 26126 18174 26178 18226
rect 26178 18174 26180 18226
rect 26124 18172 26180 18174
rect 27132 18226 27188 18228
rect 27132 18174 27134 18226
rect 27134 18174 27186 18226
rect 27186 18174 27188 18226
rect 27132 18172 27188 18174
rect 27692 17778 27748 17780
rect 27692 17726 27694 17778
rect 27694 17726 27746 17778
rect 27746 17726 27748 17778
rect 27692 17724 27748 17726
rect 24780 16828 24836 16884
rect 22764 16156 22820 16212
rect 23548 16210 23604 16212
rect 23548 16158 23550 16210
rect 23550 16158 23602 16210
rect 23602 16158 23604 16210
rect 23548 16156 23604 16158
rect 22876 15148 22932 15204
rect 24108 15148 24164 15204
rect 22092 13804 22148 13860
rect 24780 15148 24836 15204
rect 25340 17500 25396 17556
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37660 17724 37716 17780
rect 25564 16380 25620 16436
rect 26348 16828 26404 16884
rect 28140 16828 28196 16884
rect 35196 16490 35252 16492
rect 28588 16380 28644 16436
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 23212 10108 23268 10164
rect 21420 5682 21476 5684
rect 21420 5630 21422 5682
rect 21422 5630 21474 5682
rect 21474 5630 21476 5682
rect 21420 5628 21476 5630
rect 20860 4060 20916 4116
rect 22092 4114 22148 4116
rect 22092 4062 22094 4114
rect 22094 4062 22146 4114
rect 22146 4062 22148 4114
rect 22092 4060 22148 4062
rect 23772 10108 23828 10164
rect 23996 5180 24052 5236
rect 22876 3388 22932 3444
rect 24780 5234 24836 5236
rect 24780 5182 24782 5234
rect 24782 5182 24834 5234
rect 24834 5182 24836 5234
rect 24780 5180 24836 5182
rect 24892 4060 24948 4116
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 25564 3388 25620 3444
rect 25676 3612 25732 3668
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 24882 37436 24892 37492
rect 24948 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 0 36372 800 36400
rect 41200 36372 42000 36400
rect 0 36316 1708 36372
rect 1764 36316 1774 36372
rect 39778 36316 39788 36372
rect 39844 36316 42000 36372
rect 0 36288 800 36316
rect 41200 36288 42000 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 41200 35700 42000 35728
rect 40226 35644 40236 35700
rect 40292 35644 42000 35700
rect 41200 35616 42000 35644
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 20402 26908 20412 26964
rect 20468 26908 22092 26964
rect 22148 26908 22158 26964
rect 21746 26796 21756 26852
rect 21812 26796 23996 26852
rect 24052 26796 24668 26852
rect 24724 26796 25340 26852
rect 25396 26796 25406 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 0 26292 800 26320
rect 0 26236 4172 26292
rect 4228 26236 4238 26292
rect 0 26208 800 26236
rect 18162 26124 18172 26180
rect 18228 26124 19516 26180
rect 19572 26124 19582 26180
rect 23986 26124 23996 26180
rect 24052 26124 24668 26180
rect 24724 26124 24734 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 20738 25676 20748 25732
rect 20804 25676 23100 25732
rect 23156 25676 23166 25732
rect 16258 25564 16268 25620
rect 16324 25564 17500 25620
rect 17556 25564 20412 25620
rect 20468 25564 20478 25620
rect 4274 25452 4284 25508
rect 4340 25452 15372 25508
rect 15428 25452 15438 25508
rect 23426 25452 23436 25508
rect 23492 25452 24108 25508
rect 24164 25452 24174 25508
rect 16930 25340 16940 25396
rect 16996 25340 18060 25396
rect 18116 25340 18126 25396
rect 23314 25340 23324 25396
rect 23380 25340 24220 25396
rect 24276 25340 24286 25396
rect 22754 25228 22764 25284
rect 22820 25228 23772 25284
rect 23828 25228 23838 25284
rect 24098 25228 24108 25284
rect 24164 25228 25116 25284
rect 25172 25228 25182 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 0 24948 800 24976
rect 41200 24948 42000 24976
rect 0 24892 1932 24948
rect 1988 24892 1998 24948
rect 13570 24892 13580 24948
rect 13636 24892 15036 24948
rect 15092 24892 16156 24948
rect 16212 24892 16222 24948
rect 18610 24892 18620 24948
rect 18676 24892 22204 24948
rect 22260 24892 22270 24948
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 0 24864 800 24892
rect 41200 24864 42000 24892
rect 18162 24780 18172 24836
rect 18228 24780 19404 24836
rect 19460 24780 20188 24836
rect 20244 24780 20254 24836
rect 4274 24668 4284 24724
rect 4340 24668 12124 24724
rect 12180 24668 14476 24724
rect 14532 24668 15596 24724
rect 15652 24668 15662 24724
rect 19842 24668 19852 24724
rect 19908 24668 20636 24724
rect 20692 24668 20702 24724
rect 24546 24668 24556 24724
rect 24612 24668 25564 24724
rect 25620 24668 25630 24724
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 0 24192 800 24220
rect 25330 23996 25340 24052
rect 25396 23996 26796 24052
rect 26852 23996 37660 24052
rect 37716 23996 37726 24052
rect 20066 23884 20076 23940
rect 20132 23884 20412 23940
rect 20468 23884 20748 23940
rect 20804 23884 20814 23940
rect 18946 23772 18956 23828
rect 19012 23772 19628 23828
rect 19684 23772 20300 23828
rect 20356 23772 20366 23828
rect 19282 23660 19292 23716
rect 19348 23660 20188 23716
rect 20244 23660 20254 23716
rect 14130 23548 14140 23604
rect 14196 23548 19516 23604
rect 19572 23548 19582 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 19852 23324 20300 23380
rect 20356 23324 20366 23380
rect 19852 23268 19908 23324
rect 18386 23212 18396 23268
rect 18452 23212 19068 23268
rect 19124 23212 19852 23268
rect 19908 23212 19918 23268
rect 4274 23100 4284 23156
rect 4340 23100 8428 23156
rect 18498 23100 18508 23156
rect 18564 23100 19180 23156
rect 19236 23100 21308 23156
rect 21364 23100 21374 23156
rect 21634 23100 21644 23156
rect 21700 23100 22988 23156
rect 23044 23100 23054 23156
rect 23426 23100 23436 23156
rect 23492 23100 24332 23156
rect 24388 23100 24398 23156
rect 8372 23044 8428 23100
rect 8372 22988 10332 23044
rect 10388 22988 10398 23044
rect 19506 22988 19516 23044
rect 19572 22988 20188 23044
rect 20244 22988 20254 23044
rect 0 22932 800 22960
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 13458 22876 13468 22932
rect 13524 22876 14140 22932
rect 14196 22876 14206 22932
rect 14466 22876 14476 22932
rect 14532 22876 17948 22932
rect 18004 22876 18014 22932
rect 24322 22876 24332 22932
rect 24388 22876 25340 22932
rect 25396 22876 25406 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 14476 22820 14532 22876
rect 41200 22848 42000 22876
rect 12562 22764 12572 22820
rect 12628 22764 14532 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 10322 22540 10332 22596
rect 10388 22540 13468 22596
rect 13524 22540 13534 22596
rect 25554 22428 25564 22484
rect 25620 22428 26348 22484
rect 26404 22428 37660 22484
rect 37716 22428 37726 22484
rect 23538 22316 23548 22372
rect 23604 22316 25228 22372
rect 25284 22316 26796 22372
rect 26852 22316 26862 22372
rect 17938 22204 17948 22260
rect 18004 22204 20412 22260
rect 20468 22204 22092 22260
rect 22148 22204 22764 22260
rect 22820 22204 22830 22260
rect 16594 22092 16604 22148
rect 16660 22092 19516 22148
rect 19572 22092 20748 22148
rect 20804 22092 20814 22148
rect 21298 21980 21308 22036
rect 21364 21980 22204 22036
rect 22260 21980 22270 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 12786 21756 12796 21812
rect 12852 21756 13804 21812
rect 13860 21756 13870 21812
rect 18386 21756 18396 21812
rect 18452 21756 20524 21812
rect 20580 21756 20590 21812
rect 23090 21756 23100 21812
rect 23156 21756 24108 21812
rect 24164 21756 25788 21812
rect 25844 21756 25854 21812
rect 16370 21644 16380 21700
rect 16436 21644 16940 21700
rect 16996 21644 17500 21700
rect 17556 21644 19852 21700
rect 19908 21644 19918 21700
rect 20626 21644 20636 21700
rect 20692 21644 22764 21700
rect 22820 21644 22830 21700
rect 4274 21532 4284 21588
rect 4340 21532 8428 21588
rect 19618 21532 19628 21588
rect 19684 21532 22204 21588
rect 22260 21532 22270 21588
rect 26786 21532 26796 21588
rect 26852 21532 28476 21588
rect 28532 21532 37660 21588
rect 37716 21532 37726 21588
rect 8372 21476 8428 21532
rect 8372 21420 10220 21476
rect 10276 21420 10286 21476
rect 20402 21420 20412 21476
rect 20468 21420 21532 21476
rect 21588 21420 21598 21476
rect 17154 21308 17164 21364
rect 17220 21308 18396 21364
rect 18452 21308 18462 21364
rect 20962 21308 20972 21364
rect 21028 21308 22764 21364
rect 22820 21308 25564 21364
rect 25620 21308 25630 21364
rect 18834 21196 18844 21252
rect 18900 21196 20860 21252
rect 20916 21196 20926 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 20850 20972 20860 21028
rect 20916 20972 23884 21028
rect 23940 20972 23950 21028
rect 0 20916 800 20944
rect 41200 20916 42000 20944
rect 0 20860 1932 20916
rect 1988 20860 1998 20916
rect 13570 20860 13580 20916
rect 13636 20860 14924 20916
rect 14980 20860 18620 20916
rect 18676 20860 18686 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 0 20832 800 20860
rect 41200 20832 42000 20860
rect 10210 20748 10220 20804
rect 10276 20748 13468 20804
rect 13524 20748 13534 20804
rect 16034 20748 16044 20804
rect 16100 20748 17052 20804
rect 17108 20748 18508 20804
rect 18564 20748 18574 20804
rect 18946 20748 18956 20804
rect 19012 20748 20076 20804
rect 20132 20748 20142 20804
rect 17602 20636 17612 20692
rect 17668 20636 18844 20692
rect 18900 20636 18910 20692
rect 12674 20524 12684 20580
rect 12740 20524 13804 20580
rect 13860 20524 13870 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 18162 20188 18172 20244
rect 18228 20188 20412 20244
rect 20468 20188 20478 20244
rect 14802 20076 14812 20132
rect 14868 20076 15596 20132
rect 15652 20076 15662 20132
rect 20066 20076 20076 20132
rect 20132 20076 22316 20132
rect 22372 20076 22382 20132
rect 17714 19964 17724 20020
rect 17780 19964 18172 20020
rect 18228 19964 21420 20020
rect 21476 19964 23100 20020
rect 23156 19964 24108 20020
rect 24164 19964 24174 20020
rect 14018 19852 14028 19908
rect 14084 19852 15260 19908
rect 15316 19852 18060 19908
rect 18116 19852 18126 19908
rect 18386 19852 18396 19908
rect 18452 19852 21532 19908
rect 21588 19852 21868 19908
rect 21924 19852 21934 19908
rect 15810 19740 15820 19796
rect 15876 19740 16492 19796
rect 16548 19740 16558 19796
rect 21970 19740 21980 19796
rect 22036 19740 23436 19796
rect 23492 19740 26908 19796
rect 26964 19740 26974 19796
rect 15586 19628 15596 19684
rect 15652 19628 18620 19684
rect 18676 19628 23324 19684
rect 23380 19628 23390 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 4162 19292 4172 19348
rect 4228 19292 17724 19348
rect 17780 19292 18732 19348
rect 18788 19292 18798 19348
rect 24434 19292 24444 19348
rect 24500 19292 26012 19348
rect 26068 19292 26078 19348
rect 26562 19292 26572 19348
rect 26628 19292 28140 19348
rect 28196 19292 37660 19348
rect 37716 19292 37726 19348
rect 17938 19180 17948 19236
rect 18004 19180 19068 19236
rect 19124 19180 19134 19236
rect 20626 19180 20636 19236
rect 20692 19180 21756 19236
rect 21812 19180 24556 19236
rect 24612 19180 24622 19236
rect 14690 19068 14700 19124
rect 14756 19068 15820 19124
rect 15876 19068 15886 19124
rect 18946 19068 18956 19124
rect 19012 19068 22764 19124
rect 22820 19068 22830 19124
rect 12898 18956 12908 19012
rect 12964 18956 13692 19012
rect 13748 18956 13758 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 18050 18508 18060 18564
rect 18116 18508 18564 18564
rect 24546 18508 24556 18564
rect 24612 18508 25900 18564
rect 25956 18508 25966 18564
rect 18508 18452 18564 18508
rect 11554 18396 11564 18452
rect 11620 18396 14028 18452
rect 14084 18396 14812 18452
rect 14868 18396 15484 18452
rect 15540 18396 15550 18452
rect 18508 18396 19404 18452
rect 19460 18396 19470 18452
rect 23874 18396 23884 18452
rect 23940 18396 25340 18452
rect 25396 18396 25406 18452
rect 14354 18284 14364 18340
rect 14420 18284 16044 18340
rect 16100 18284 16110 18340
rect 16818 18284 16828 18340
rect 16884 18284 18060 18340
rect 18116 18284 18126 18340
rect 19282 18284 19292 18340
rect 19348 18284 19964 18340
rect 20020 18284 20972 18340
rect 21028 18284 21038 18340
rect 24658 18284 24668 18340
rect 24724 18284 26348 18340
rect 26404 18284 26414 18340
rect 41200 18228 42000 18256
rect 14914 18172 14924 18228
rect 14980 18172 16268 18228
rect 16324 18172 20860 18228
rect 20916 18172 22092 18228
rect 22148 18172 25564 18228
rect 25620 18172 25630 18228
rect 26114 18172 26124 18228
rect 26180 18172 27132 18228
rect 27188 18172 27198 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19394 17836 19404 17892
rect 19460 17836 21644 17892
rect 21700 17836 21710 17892
rect 1922 17724 1932 17780
rect 1988 17724 1998 17780
rect 27682 17724 27692 17780
rect 27748 17724 37660 17780
rect 37716 17724 37726 17780
rect 0 17556 800 17584
rect 1932 17556 1988 17724
rect 4274 17612 4284 17668
rect 4340 17612 12460 17668
rect 12516 17612 15596 17668
rect 15652 17612 15662 17668
rect 16370 17612 16380 17668
rect 16436 17612 19852 17668
rect 19908 17612 19918 17668
rect 20132 17612 20636 17668
rect 20692 17612 21868 17668
rect 21924 17612 21934 17668
rect 20132 17556 20188 17612
rect 0 17500 1988 17556
rect 14242 17500 14252 17556
rect 14308 17500 15372 17556
rect 15428 17500 20188 17556
rect 22194 17500 22204 17556
rect 22260 17500 25340 17556
rect 25396 17500 25406 17556
rect 0 17472 800 17500
rect 14578 17388 14588 17444
rect 14644 17388 16268 17444
rect 16324 17388 16334 17444
rect 19954 17388 19964 17444
rect 20020 17388 20748 17444
rect 20804 17388 20814 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 15698 17164 15708 17220
rect 15764 17164 17612 17220
rect 17668 17164 18732 17220
rect 18788 17164 18798 17220
rect 20738 17164 20748 17220
rect 20804 17164 21420 17220
rect 21476 17164 21486 17220
rect 16482 17052 16492 17108
rect 16548 17052 17276 17108
rect 17332 17052 17342 17108
rect 19506 17052 19516 17108
rect 19572 17052 19908 17108
rect 20402 17052 20412 17108
rect 20468 17052 22092 17108
rect 22148 17052 23100 17108
rect 23156 17052 23166 17108
rect 14690 16940 14700 16996
rect 14756 16940 16604 16996
rect 16660 16940 16670 16996
rect 19852 16884 19908 17052
rect 20066 16940 20076 16996
rect 20132 16940 20748 16996
rect 20804 16940 20814 16996
rect 15810 16828 15820 16884
rect 15876 16828 17500 16884
rect 17556 16828 17566 16884
rect 18610 16828 18620 16884
rect 18676 16828 19628 16884
rect 19684 16828 19694 16884
rect 19852 16828 20300 16884
rect 20356 16828 22428 16884
rect 22484 16828 22494 16884
rect 24770 16828 24780 16884
rect 24836 16828 26348 16884
rect 26404 16828 28140 16884
rect 28196 16828 28206 16884
rect 18498 16716 18508 16772
rect 18564 16716 19180 16772
rect 19236 16716 20524 16772
rect 20580 16716 20590 16772
rect 20066 16604 20076 16660
rect 20132 16604 21420 16660
rect 21476 16604 21486 16660
rect 20710 16492 20748 16548
rect 20804 16492 20814 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 25554 16380 25564 16436
rect 25620 16380 28588 16436
rect 28644 16380 28654 16436
rect 22754 16156 22764 16212
rect 22820 16156 23548 16212
rect 23604 16156 23614 16212
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 20626 15372 20636 15428
rect 20692 15372 21532 15428
rect 21588 15372 21598 15428
rect 19506 15148 19516 15204
rect 19572 15148 20188 15204
rect 20244 15148 20254 15204
rect 20850 15148 20860 15204
rect 20916 15148 22876 15204
rect 22932 15148 24108 15204
rect 24164 15148 24780 15204
rect 24836 15148 24846 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 14690 14252 14700 14308
rect 14756 14252 16380 14308
rect 16436 14252 16446 14308
rect 18274 14252 18284 14308
rect 18340 14252 19404 14308
rect 19460 14252 19470 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 17378 13804 17388 13860
rect 17444 13804 22092 13860
rect 22148 13804 22158 13860
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 16482 13132 16492 13188
rect 16548 13132 17164 13188
rect 17220 13132 17230 13188
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 23202 10108 23212 10164
rect 23268 10108 23772 10164
rect 23828 10108 23838 10164
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 20178 5628 20188 5684
rect 20244 5628 21420 5684
rect 21476 5628 21486 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 16818 5180 16828 5236
rect 16884 5180 18060 5236
rect 18116 5180 18126 5236
rect 23986 5180 23996 5236
rect 24052 5180 24780 5236
rect 24836 5180 24846 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 17714 4060 17724 4116
rect 17780 4060 18732 4116
rect 18788 4060 18798 4116
rect 20850 4060 20860 4116
rect 20916 4060 22092 4116
rect 22148 4060 22158 4116
rect 24882 4060 24892 4116
rect 24948 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 25666 3612 25676 3668
rect 25732 3612 29372 3668
rect 29428 3612 29438 3668
rect 22866 3388 22876 3444
rect 22932 3388 25564 3444
rect 25620 3388 25630 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 20748 16940 20804 16996
rect 20748 16492 20804 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 20748 16996 20804 17006
rect 20748 16548 20804 16940
rect 20748 16482 20804 16492
rect 35168 16492 35488 18004
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _082_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18592 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _083_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _084_
timestamp 1698175906
transform 1 0 16016 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _085_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16800 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _086_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16128 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _087_
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _088_
timestamp 1698175906
transform -1 0 15120 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _089_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _090_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13104 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _091_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _092_
timestamp 1698175906
transform 1 0 19040 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _093_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20048 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _095_
timestamp 1698175906
transform 1 0 18032 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19712 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _097_
timestamp 1698175906
transform 1 0 13440 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _098_
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform -1 0 20384 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18256 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _101_
timestamp 1698175906
transform 1 0 17696 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _102_
timestamp 1698175906
transform -1 0 13104 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21280 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19936 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _105_
timestamp 1698175906
transform -1 0 19712 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _106_
timestamp 1698175906
transform -1 0 23632 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _107_
timestamp 1698175906
transform -1 0 20944 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform 1 0 20048 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _109_
timestamp 1698175906
transform 1 0 21840 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22400 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_
timestamp 1698175906
transform 1 0 21504 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _112_
timestamp 1698175906
transform 1 0 22736 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _113_
timestamp 1698175906
transform 1 0 22400 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _114_
timestamp 1698175906
transform 1 0 13328 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _115_
timestamp 1698175906
transform -1 0 12992 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _116_
timestamp 1698175906
transform 1 0 22736 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _117_
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_
timestamp 1698175906
transform -1 0 24752 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _119_
timestamp 1698175906
transform -1 0 15008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13776 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _121_
timestamp 1698175906
transform 1 0 26880 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _122_
timestamp 1698175906
transform -1 0 26320 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_
timestamp 1698175906
transform -1 0 26880 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _124_
timestamp 1698175906
transform -1 0 24864 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform -1 0 27104 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _126_
timestamp 1698175906
transform 1 0 25424 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _127_
timestamp 1698175906
transform -1 0 20384 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _128_
timestamp 1698175906
transform -1 0 17584 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698175906
transform -1 0 16688 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1698175906
transform -1 0 17808 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17808 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _132_
timestamp 1698175906
transform -1 0 16912 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _133_
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _134_
timestamp 1698175906
transform -1 0 22064 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21168 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _136_
timestamp 1698175906
transform -1 0 20832 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform 1 0 20160 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 22624 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _140_
timestamp 1698175906
transform 1 0 16128 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _141_
timestamp 1698175906
transform -1 0 18704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 20384 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _143_
timestamp 1698175906
transform 1 0 18256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _145_
timestamp 1698175906
transform 1 0 22848 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _147_
timestamp 1698175906
transform 1 0 23744 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 24304 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20048 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21840 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform 1 0 22512 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform -1 0 22400 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _153_
timestamp 1698175906
transform -1 0 21504 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698175906
transform 1 0 19824 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform 1 0 16800 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform -1 0 19376 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _158_
timestamp 1698175906
transform -1 0 19040 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _159_
timestamp 1698175906
transform 1 0 19376 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform -1 0 20160 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _163_
timestamp 1698175906
transform -1 0 22512 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23296 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _165_
timestamp 1698175906
transform 1 0 21616 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _166_
timestamp 1698175906
transform -1 0 15568 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _167_
timestamp 1698175906
transform 1 0 13888 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _168_
timestamp 1698175906
transform 1 0 11312 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _169_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _170_
timestamp 1698175906
transform 1 0 16016 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _171_
timestamp 1698175906
transform -1 0 13328 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _172_
timestamp 1698175906
transform 1 0 17360 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _173_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22624 0 1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _175_
timestamp 1698175906
transform -1 0 13440 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _176_
timestamp 1698175906
transform 1 0 23744 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _177_
timestamp 1698175906
transform -1 0 15232 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _178_
timestamp 1698175906
transform 1 0 24640 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _179_
timestamp 1698175906
transform 1 0 25088 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _180_
timestamp 1698175906
transform 1 0 25424 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _181_
timestamp 1698175906
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_
timestamp 1698175906
transform 1 0 13776 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1698175906
transform 1 0 20608 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1698175906
transform 1 0 17696 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _189_
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _190_
timestamp 1698175906
transform -1 0 15904 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _191_
timestamp 1698175906
transform 1 0 17024 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _192_
timestamp 1698175906
transform 1 0 22736 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _193_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__CLK
timestamp 1698175906
transform 1 0 15792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__CLK
timestamp 1698175906
transform 1 0 17360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__CLK
timestamp 1698175906
transform -1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__CLK
timestamp 1698175906
transform 1 0 20384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__CLK
timestamp 1698175906
transform -1 0 18032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__CLK
timestamp 1698175906
transform 1 0 24640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__CLK
timestamp 1698175906
transform 1 0 26320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__CLK
timestamp 1698175906
transform 1 0 13552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__CLK
timestamp 1698175906
transform 1 0 27216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__CLK
timestamp 1698175906
transform 1 0 16128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__CLK
timestamp 1698175906
transform 1 0 28112 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__CLK
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__CLK
timestamp 1698175906
transform 1 0 28896 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__CLK
timestamp 1698175906
transform 1 0 17920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__CLK
timestamp 1698175906
transform 1 0 24080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK
timestamp 1698175906
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 17808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18592 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20720 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22176 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698175906
transform 1 0 31136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698175906
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698175906
transform 1 0 17472 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_171
timestamp 1698175906
transform 1 0 20496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_201 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23856 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_165
timestamp 1698175906
transform 1 0 19824 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_173
timestamp 1698175906
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698175906
transform 1 0 22960 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_197
timestamp 1698175906
transform 1 0 23408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_225
timestamp 1698175906
transform 1 0 26544 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_158
timestamp 1698175906
transform 1 0 19040 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_166
timestamp 1698175906
transform 1 0 19936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_168
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_195
timestamp 1698175906
transform 1 0 23184 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_203
timestamp 1698175906
transform 1 0 24080 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_207
timestamp 1698175906
transform 1 0 24528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698175906
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_145
timestamp 1698175906
transform 1 0 17584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_149
timestamp 1698175906
transform 1 0 18032 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_165
timestamp 1698175906
transform 1 0 19824 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_185
timestamp 1698175906
transform 1 0 22064 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_189
timestamp 1698175906
transform 1 0 22512 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_197
timestamp 1698175906
transform 1 0 23408 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_229
timestamp 1698175906
transform 1 0 26992 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_201
timestamp 1698175906
transform 1 0 23856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_205
timestamp 1698175906
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_137
timestamp 1698175906
transform 1 0 16688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_139
timestamp 1698175906
transform 1 0 16912 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_146
timestamp 1698175906
transform 1 0 17696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_150
timestamp 1698175906
transform 1 0 18144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_164
timestamp 1698175906
transform 1 0 19712 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_191
timestamp 1698175906
transform 1 0 22736 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_223
timestamp 1698175906
transform 1 0 26320 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_162
timestamp 1698175906
transform 1 0 19488 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_180
timestamp 1698175906
transform 1 0 21504 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_196
timestamp 1698175906
transform 1 0 23296 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698175906
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_218
timestamp 1698175906
transform 1 0 25760 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_250
timestamp 1698175906
transform 1 0 29344 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_266
timestamp 1698175906
transform 1 0 31136 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698175906
transform 1 0 32032 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_140
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_189
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_221
timestamp 1698175906
transform 1 0 26096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_225
timestamp 1698175906
transform 1 0 26544 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_96
timestamp 1698175906
transform 1 0 12096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_127
timestamp 1698175906
transform 1 0 15568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_147
timestamp 1698175906
transform 1 0 17808 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_163
timestamp 1698175906
transform 1 0 19600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_177
timestamp 1698175906
transform 1 0 21168 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_181
timestamp 1698175906
transform 1 0 21616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_188
timestamp 1698175906
transform 1 0 22400 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_204
timestamp 1698175906
transform 1 0 24192 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_218
timestamp 1698175906
transform 1 0 25760 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_250
timestamp 1698175906
transform 1 0 29344 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_266
timestamp 1698175906
transform 1 0 31136 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698175906
transform 1 0 32032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698175906
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_121
timestamp 1698175906
transform 1 0 14896 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_137
timestamp 1698175906
transform 1 0 16688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_145
timestamp 1698175906
transform 1 0 17584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_149
timestamp 1698175906
transform 1 0 18032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_158
timestamp 1698175906
transform 1 0 19040 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_162
timestamp 1698175906
transform 1 0 19488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_196
timestamp 1698175906
transform 1 0 23296 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_204
timestamp 1698175906
transform 1 0 24192 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_237
timestamp 1698175906
transform 1 0 27888 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_118
timestamp 1698175906
transform 1 0 14560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_122
timestamp 1698175906
transform 1 0 15008 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_126
timestamp 1698175906
transform 1 0 15456 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_128
timestamp 1698175906
transform 1 0 15680 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_178
timestamp 1698175906
transform 1 0 21280 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_233
timestamp 1698175906
transform 1 0 27440 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_265
timestamp 1698175906
transform 1 0 31024 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698175906
transform 1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698175906
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_93
timestamp 1698175906
transform 1 0 11760 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_97
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_188
timestamp 1698175906
transform 1 0 22400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_190
timestamp 1698175906
transform 1 0 22624 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_210
timestamp 1698175906
transform 1 0 24864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_241
timestamp 1698175906
transform 1 0 28336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_120
timestamp 1698175906
transform 1 0 14784 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_124
timestamp 1698175906
transform 1 0 15232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_132
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_204
timestamp 1698175906
transform 1 0 24192 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_244
timestamp 1698175906
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_248
timestamp 1698175906
transform 1 0 29120 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698175906
transform 1 0 9072 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_85
timestamp 1698175906
transform 1 0 10864 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_93
timestamp 1698175906
transform 1 0 11760 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_97
timestamp 1698175906
transform 1 0 12208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_116
timestamp 1698175906
transform 1 0 14336 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_179
timestamp 1698175906
transform 1 0 21392 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_236
timestamp 1698175906
transform 1 0 27776 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698175906
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_76
timestamp 1698175906
transform 1 0 9856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_116
timestamp 1698175906
transform 1 0 14336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_120
timestamp 1698175906
transform 1 0 14784 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_189
timestamp 1698175906
transform 1 0 22512 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_198
timestamp 1698175906
transform 1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698175906
transform 1 0 25312 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_223
timestamp 1698175906
transform 1 0 26320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_230
timestamp 1698175906
transform 1 0 27104 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_262
timestamp 1698175906
transform 1 0 30688 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_85
timestamp 1698175906
transform 1 0 10864 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_93
timestamp 1698175906
transform 1 0 11760 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_97
timestamp 1698175906
transform 1 0 12208 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698175906
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_141
timestamp 1698175906
transform 1 0 17136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_145
timestamp 1698175906
transform 1 0 17584 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_155
timestamp 1698175906
transform 1 0 18704 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_159
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698175906
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_188
timestamp 1698175906
transform 1 0 22400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_225
timestamp 1698175906
transform 1 0 26544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_229
timestamp 1698175906
transform 1 0 26992 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_76
timestamp 1698175906
transform 1 0 9856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_78
timestamp 1698175906
transform 1 0 10080 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_108
timestamp 1698175906
transform 1 0 13440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_110
timestamp 1698175906
transform 1 0 13664 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_121
timestamp 1698175906
transform 1 0 14896 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_150
timestamp 1698175906
transform 1 0 18144 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_161
timestamp 1698175906
transform 1 0 19376 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_178
timestamp 1698175906
transform 1 0 21280 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_186
timestamp 1698175906
transform 1 0 22176 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_190
timestamp 1698175906
transform 1 0 22624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_198
timestamp 1698175906
transform 1 0 23520 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698175906
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_217
timestamp 1698175906
transform 1 0 25648 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_249
timestamp 1698175906
transform 1 0 29232 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_265
timestamp 1698175906
transform 1 0 31024 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_111
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_122
timestamp 1698175906
transform 1 0 15008 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_154
timestamp 1698175906
transform 1 0 18592 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_164
timestamp 1698175906
transform 1 0 19712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_193
timestamp 1698175906
transform 1 0 22960 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_197
timestamp 1698175906
transform 1 0 23408 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_199
timestamp 1698175906
transform 1 0 23632 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_229
timestamp 1698175906
transform 1 0 26992 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_233
timestamp 1698175906
transform 1 0 27440 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 11200 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_92
timestamp 1698175906
transform 1 0 11648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_94
timestamp 1698175906
transform 1 0 11872 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_130
timestamp 1698175906
transform 1 0 15904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698175906
transform 1 0 16352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_146
timestamp 1698175906
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_148
timestamp 1698175906
transform 1 0 17920 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_157
timestamp 1698175906
transform 1 0 18928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_172
timestamp 1698175906
transform 1 0 20608 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_217
timestamp 1698175906
transform 1 0 25648 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_249
timestamp 1698175906
transform 1 0 29232 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_265
timestamp 1698175906
transform 1 0 31024 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 31920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_123
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_168
timestamp 1698175906
transform 1 0 20160 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 22064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_199
timestamp 1698175906
transform 1 0 23632 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_205
timestamp 1698175906
transform 1 0 24304 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_237
timestamp 1698175906
transform 1 0 27888 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_136
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_179
timestamp 1698175906
transform 1 0 21392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_216
timestamp 1698175906
transform 1 0 25536 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_139
timestamp 1698175906
transform 1 0 16912 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_155
timestamp 1698175906
transform 1 0 18704 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_163
timestamp 1698175906
transform 1 0 19600 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_167
timestamp 1698175906
transform 1 0 20048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_169
timestamp 1698175906
transform 1 0 20272 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_206
timestamp 1698175906
transform 1 0 24416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_210
timestamp 1698175906
transform 1 0 24864 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698175906
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698175906
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698175906
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698175906
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698175906
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita45_23 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita45_24
timestamp 1698175906
transform 1 0 20832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita45_25
timestamp 1698175906
transform 1 0 39984 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita45_26
timestamp 1698175906
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16912 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 23632 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 24192 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 20944 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 17584 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 20272 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 4480 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 41200 36288 42000 36400 0 FreeSans 448 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 41200 35616 42000 35728 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 24024 22008 24024 22008 0 _000_
rlabel metal2 22792 25928 22792 25928 0 _001_
rlabel metal2 14616 17192 14616 17192 0 _002_
rlabel metal2 23352 20664 23352 20664 0 _003_
rlabel metal2 12264 18760 12264 18760 0 _004_
rlabel metal2 19544 25872 19544 25872 0 _005_
rlabel metal2 18312 25144 18312 25144 0 _006_
rlabel metal2 12600 21224 12600 21224 0 _007_
rlabel metal2 18312 14056 18312 14056 0 _008_
rlabel metal3 21280 26936 21280 26936 0 _009_
rlabel metal3 23184 16184 23184 16184 0 _010_
rlabel metal2 12488 22792 12488 22792 0 _011_
rlabel metal2 24696 24248 24696 24248 0 _012_
rlabel metal2 14280 23968 14280 23968 0 _013_
rlabel metal2 25648 17752 25648 17752 0 _014_
rlabel metal3 25256 19320 25256 19320 0 _015_
rlabel metal2 25704 20804 25704 20804 0 _016_
rlabel metal2 14728 14056 14728 14056 0 _017_
rlabel metal2 14728 16576 14728 16576 0 _018_
rlabel metal2 21560 14056 21560 14056 0 _019_
rlabel metal2 19768 17416 19768 17416 0 _020_
rlabel metal2 23016 18312 23016 18312 0 _021_
rlabel metal3 13328 21784 13328 21784 0 _022_
rlabel metal2 23464 22456 23464 22456 0 _023_
rlabel metal3 25088 24696 25088 24696 0 _024_
rlabel metal2 14728 23408 14728 23408 0 _025_
rlabel metal3 26656 18200 26656 18200 0 _026_
rlabel metal2 26376 18368 26376 18368 0 _027_
rlabel metal2 26432 21560 26432 21560 0 _028_
rlabel metal3 19880 16968 19880 16968 0 _029_
rlabel metal2 17192 13104 17192 13104 0 _030_
rlabel metal3 16912 17080 16912 17080 0 _031_
rlabel metal2 16856 17584 16856 17584 0 _032_
rlabel metal2 21896 14560 21896 14560 0 _033_
rlabel metal2 20216 17360 20216 17360 0 _034_
rlabel metal2 20440 23520 20440 23520 0 _035_
rlabel metal2 20440 22568 20440 22568 0 _036_
rlabel metal3 23632 21784 23632 21784 0 _037_
rlabel metal2 20776 22736 20776 22736 0 _038_
rlabel metal2 20552 21280 20552 21280 0 _039_
rlabel metal2 20888 20888 20888 20888 0 _040_
rlabel metal2 21336 22848 21336 22848 0 _041_
rlabel metal2 21672 22848 21672 22848 0 _042_
rlabel metal2 25256 23968 25256 23968 0 _043_
rlabel metal2 24360 22344 24360 22344 0 _044_
rlabel metal3 23296 25256 23296 25256 0 _045_
rlabel metal2 20216 21168 20216 21168 0 _046_
rlabel metal2 22232 23856 22232 23856 0 _047_
rlabel metal2 21840 22120 21840 22120 0 _048_
rlabel metal2 20944 15512 20944 15512 0 _049_
rlabel metal2 18984 23464 18984 23464 0 _050_
rlabel metal2 20888 22176 20888 22176 0 _051_
rlabel metal3 21896 21336 21896 21336 0 _052_
rlabel metal2 18872 23408 18872 23408 0 _053_
rlabel metal2 17640 17080 17640 17080 0 _054_
rlabel metal2 20216 21952 20216 21952 0 _055_
rlabel metal2 21448 19600 21448 19600 0 _056_
rlabel metal2 21952 16968 21952 16968 0 _057_
rlabel metal2 19600 20776 19600 20776 0 _058_
rlabel metal2 21952 21672 21952 21672 0 _059_
rlabel metal3 16072 19880 16072 19880 0 _060_
rlabel metal2 15960 17752 15960 17752 0 _061_
rlabel metal2 15848 19544 15848 19544 0 _062_
rlabel metal2 22008 17920 22008 17920 0 _063_
rlabel metal2 13944 21168 13944 21168 0 _064_
rlabel metal2 12936 19040 12936 19040 0 _065_
rlabel metal2 18032 21336 18032 21336 0 _066_
rlabel metal2 20216 23856 20216 23856 0 _067_
rlabel metal2 20664 25928 20664 25928 0 _068_
rlabel metal2 13608 21560 13608 21560 0 _069_
rlabel metal2 13720 21952 13720 21952 0 _070_
rlabel metal3 13272 20552 13272 20552 0 _071_
rlabel metal2 19768 20552 19768 20552 0 _072_
rlabel metal2 17864 21560 17864 21560 0 _073_
rlabel metal3 16240 22904 16240 22904 0 _074_
rlabel metal2 20664 16184 20664 16184 0 _075_
rlabel metal3 19880 15176 19880 15176 0 _076_
rlabel metal2 23128 25592 23128 25592 0 _077_
rlabel metal2 22792 21616 22792 21616 0 _078_
rlabel metal2 22344 17136 22344 17136 0 _079_
rlabel metal2 22120 17808 22120 17808 0 _080_
rlabel metal2 23464 19488 23464 19488 0 _081_
rlabel metal3 2478 26264 2478 26264 0 clk
rlabel metal2 22344 20440 22344 20440 0 clknet_0_clk
rlabel metal2 17528 25928 17528 25928 0 clknet_1_0__leaf_clk
rlabel metal2 21840 26264 21840 26264 0 clknet_1_1__leaf_clk
rlabel metal2 17528 21616 17528 21616 0 dut45.count\[0\]
rlabel metal2 18536 21896 18536 21896 0 dut45.count\[1\]
rlabel metal2 20664 24304 20664 24304 0 dut45.count\[2\]
rlabel metal2 20328 23324 20328 23324 0 dut45.count\[3\]
rlabel metal2 17472 17080 17472 17080 0 net1
rlabel metal2 17248 12824 17248 12824 0 net10
rlabel metal2 25368 24416 25368 24416 0 net11
rlabel metal2 26600 18984 26600 18984 0 net12
rlabel metal2 26824 21616 26824 21616 0 net13
rlabel metal3 6356 23128 6356 23128 0 net14
rlabel metal3 27104 16408 27104 16408 0 net15
rlabel metal3 23800 25368 23800 25368 0 net16
rlabel metal2 20440 9744 20440 9744 0 net17
rlabel metal3 6356 21560 6356 21560 0 net18
rlabel metal2 12488 17192 12488 17192 0 net19
rlabel metal2 23240 11424 23240 11424 0 net2
rlabel metal2 24752 26152 24752 26152 0 net20
rlabel metal2 27216 18536 27216 18536 0 net21
rlabel metal2 25424 23240 25424 23240 0 net22
rlabel metal3 40530 36344 40530 36344 0 net23
rlabel metal2 21560 2030 21560 2030 0 net24
rlabel metal2 40264 35952 40264 35952 0 net25
rlabel metal3 1246 36344 1246 36344 0 net26
rlabel metal2 23352 12936 23352 12936 0 net3
rlabel metal4 20776 16744 20776 16744 0 net4
rlabel metal2 25592 9856 25592 9856 0 net5
rlabel metal2 25816 15736 25816 15736 0 net6
rlabel metal2 15400 25200 15400 25200 0 net7
rlabel metal2 12152 24640 12152 24640 0 net8
rlabel metal2 17528 8904 17528 8904 0 net9
rlabel metal3 17472 5208 17472 5208 0 segm[10]
rlabel metal2 23576 854 23576 854 0 segm[11]
rlabel metal2 22232 2086 22232 2086 0 segm[12]
rlabel metal3 21504 4088 21504 4088 0 segm[13]
rlabel metal3 25592 4088 25592 4088 0 segm[3]
rlabel metal3 24248 3416 24248 3416 0 segm[5]
rlabel metal3 1358 24920 1358 24920 0 segm[6]
rlabel metal3 1358 24248 1358 24248 0 segm[7]
rlabel metal2 18200 2058 18200 2058 0 segm[8]
rlabel metal2 17528 2058 17528 2058 0 segm[9]
rlabel metal2 40040 25256 40040 25256 0 sel[0]
rlabel metal2 40040 19656 40040 19656 0 sel[10]
rlabel metal2 40040 21112 40040 21112 0 sel[11]
rlabel metal3 1358 22904 1358 22904 0 sel[1]
rlabel metal2 25592 1190 25592 1190 0 sel[2]
rlabel metal2 22904 39746 22904 39746 0 sel[3]
rlabel metal3 20832 5656 20832 5656 0 sel[4]
rlabel metal3 1358 20888 1358 20888 0 sel[5]
rlabel metal3 1358 17528 1358 17528 0 sel[6]
rlabel metal2 24920 39354 24920 39354 0 sel[7]
rlabel metal3 40642 18200 40642 18200 0 sel[8]
rlabel metal3 40642 22904 40642 22904 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
