magic
tech gf180mcuD
magscale 1 10
timestamp 1699643791
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 15374 38274 15426 38286
rect 15374 38210 15426 38222
rect 19182 38274 19234 38286
rect 19182 38210 19234 38222
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 15922 37998 15934 38050
rect 15986 37998 15998 38050
rect 19730 37998 19742 38050
rect 19794 37998 19806 38050
rect 21410 37998 21422 38050
rect 21474 37998 21486 38050
rect 24994 37998 25006 38050
rect 25058 37998 25070 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 22766 37490 22818 37502
rect 22766 37426 22818 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 21186 37214 21198 37266
rect 21250 37214 21262 37266
rect 21858 37214 21870 37266
rect 21922 37214 21934 37266
rect 25554 37214 25566 37266
rect 25618 37214 25630 37266
rect 20066 37102 20078 37154
rect 20130 37102 20142 37154
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 18062 36706 18114 36718
rect 18062 36642 18114 36654
rect 22318 36706 22370 36718
rect 22318 36642 22370 36654
rect 26126 36706 26178 36718
rect 26126 36642 26178 36654
rect 17154 36430 17166 36482
rect 17218 36430 17230 36482
rect 21746 36430 21758 36482
rect 21810 36430 21822 36482
rect 25218 36430 25230 36482
rect 25282 36430 25294 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 14478 28418 14530 28430
rect 14478 28354 14530 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 14814 28082 14866 28094
rect 14814 28018 14866 28030
rect 15598 27858 15650 27870
rect 14130 27806 14142 27858
rect 14194 27806 14206 27858
rect 15026 27806 15038 27858
rect 15090 27806 15102 27858
rect 15362 27806 15374 27858
rect 15426 27806 15438 27858
rect 15598 27794 15650 27806
rect 16046 27858 16098 27870
rect 22318 27858 22370 27870
rect 18946 27806 18958 27858
rect 19010 27806 19022 27858
rect 16046 27794 16098 27806
rect 22318 27794 22370 27806
rect 17502 27746 17554 27758
rect 11218 27694 11230 27746
rect 11282 27694 11294 27746
rect 13346 27694 13358 27746
rect 13410 27694 13422 27746
rect 19618 27694 19630 27746
rect 19682 27694 19694 27746
rect 21746 27694 21758 27746
rect 21810 27694 21822 27746
rect 17502 27682 17554 27694
rect 15150 27634 15202 27646
rect 15150 27570 15202 27582
rect 15934 27634 15986 27646
rect 15934 27570 15986 27582
rect 16046 27634 16098 27646
rect 16046 27570 16098 27582
rect 16494 27634 16546 27646
rect 16494 27570 16546 27582
rect 16718 27634 16770 27646
rect 16718 27570 16770 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 1934 27186 1986 27198
rect 25006 27186 25058 27198
rect 15026 27134 15038 27186
rect 15090 27134 15102 27186
rect 17154 27134 17166 27186
rect 17218 27134 17230 27186
rect 20514 27134 20526 27186
rect 20578 27134 20590 27186
rect 1934 27122 1986 27134
rect 25006 27122 25058 27134
rect 25678 27074 25730 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 14242 27022 14254 27074
rect 14306 27022 14318 27074
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 22194 27022 22206 27074
rect 22258 27022 22270 27074
rect 25678 27010 25730 27022
rect 21310 26962 21362 26974
rect 18386 26910 18398 26962
rect 18450 26910 18462 26962
rect 21310 26898 21362 26910
rect 21422 26962 21474 26974
rect 21422 26898 21474 26910
rect 21646 26962 21698 26974
rect 22866 26910 22878 26962
rect 22930 26910 22942 26962
rect 21646 26898 21698 26910
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 16158 26514 16210 26526
rect 16158 26450 16210 26462
rect 16270 26514 16322 26526
rect 16270 26450 16322 26462
rect 18734 26514 18786 26526
rect 18734 26450 18786 26462
rect 19742 26514 19794 26526
rect 19742 26450 19794 26462
rect 20750 26514 20802 26526
rect 20750 26450 20802 26462
rect 22318 26514 22370 26526
rect 22318 26450 22370 26462
rect 23662 26514 23714 26526
rect 23662 26450 23714 26462
rect 24334 26514 24386 26526
rect 25230 26514 25282 26526
rect 24658 26462 24670 26514
rect 24722 26462 24734 26514
rect 25554 26462 25566 26514
rect 25618 26462 25630 26514
rect 24334 26450 24386 26462
rect 25230 26450 25282 26462
rect 19518 26402 19570 26414
rect 13794 26350 13806 26402
rect 13858 26350 13870 26402
rect 19518 26338 19570 26350
rect 19966 26402 20018 26414
rect 19966 26338 20018 26350
rect 21310 26402 21362 26414
rect 22430 26402 22482 26414
rect 21634 26350 21646 26402
rect 21698 26350 21710 26402
rect 21310 26338 21362 26350
rect 22430 26338 22482 26350
rect 16830 26290 16882 26302
rect 13122 26238 13134 26290
rect 13186 26238 13198 26290
rect 16482 26238 16494 26290
rect 16546 26238 16558 26290
rect 16830 26226 16882 26238
rect 18510 26290 18562 26302
rect 18510 26226 18562 26238
rect 18846 26290 18898 26302
rect 18846 26226 18898 26238
rect 19182 26290 19234 26302
rect 19182 26226 19234 26238
rect 20414 26290 20466 26302
rect 20414 26226 20466 26238
rect 20750 26290 20802 26302
rect 20750 26226 20802 26238
rect 21086 26290 21138 26302
rect 21086 26226 21138 26238
rect 22206 26290 22258 26302
rect 22206 26226 22258 26238
rect 22878 26290 22930 26302
rect 22878 26226 22930 26238
rect 23438 26290 23490 26302
rect 23438 26226 23490 26238
rect 23774 26290 23826 26302
rect 23774 26226 23826 26238
rect 17502 26178 17554 26190
rect 15922 26126 15934 26178
rect 15986 26126 15998 26178
rect 17502 26114 17554 26126
rect 19630 26178 19682 26190
rect 19630 26114 19682 26126
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 14814 25730 14866 25742
rect 14814 25666 14866 25678
rect 15710 25730 15762 25742
rect 15710 25666 15762 25678
rect 15822 25618 15874 25630
rect 15822 25554 15874 25566
rect 14142 25394 14194 25406
rect 14142 25330 14194 25342
rect 14254 25394 14306 25406
rect 14254 25330 14306 25342
rect 14478 25394 14530 25406
rect 14478 25330 14530 25342
rect 14702 25394 14754 25406
rect 14702 25330 14754 25342
rect 15150 25394 15202 25406
rect 19842 25342 19854 25394
rect 19906 25342 19918 25394
rect 15150 25330 15202 25342
rect 14926 25282 14978 25294
rect 14926 25218 14978 25230
rect 16270 25282 16322 25294
rect 16270 25218 16322 25230
rect 20190 25282 20242 25294
rect 20190 25218 20242 25230
rect 20638 25282 20690 25294
rect 20638 25218 20690 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 17614 24946 17666 24958
rect 17614 24882 17666 24894
rect 20750 24946 20802 24958
rect 21074 24894 21086 24946
rect 21138 24894 21150 24946
rect 20750 24882 20802 24894
rect 14366 24722 14418 24734
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 14366 24658 14418 24670
rect 10994 24558 11006 24610
rect 11058 24558 11070 24610
rect 13122 24558 13134 24610
rect 13186 24558 13198 24610
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 1934 24050 1986 24062
rect 1934 23986 1986 23998
rect 15934 24050 15986 24062
rect 15934 23986 15986 23998
rect 19518 24050 19570 24062
rect 40014 24050 40066 24062
rect 26114 23998 26126 24050
rect 26178 23998 26190 24050
rect 19518 23986 19570 23998
rect 40014 23986 40066 23998
rect 15486 23938 15538 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 15486 23874 15538 23886
rect 16158 23938 16210 23950
rect 16706 23886 16718 23938
rect 16770 23886 16782 23938
rect 21410 23886 21422 23938
rect 21474 23886 21486 23938
rect 23202 23886 23214 23938
rect 23266 23886 23278 23938
rect 37874 23886 37886 23938
rect 37938 23886 37950 23938
rect 16158 23874 16210 23886
rect 14366 23826 14418 23838
rect 14366 23762 14418 23774
rect 14478 23826 14530 23838
rect 14478 23762 14530 23774
rect 15710 23826 15762 23838
rect 15710 23762 15762 23774
rect 17278 23826 17330 23838
rect 17278 23762 17330 23774
rect 19406 23826 19458 23838
rect 21634 23774 21646 23826
rect 21698 23774 21710 23826
rect 23986 23774 23998 23826
rect 24050 23774 24062 23826
rect 19406 23762 19458 23774
rect 14142 23714 14194 23726
rect 14142 23650 14194 23662
rect 15598 23714 15650 23726
rect 19630 23714 19682 23726
rect 16482 23662 16494 23714
rect 16546 23662 16558 23714
rect 15598 23650 15650 23662
rect 19630 23650 19682 23662
rect 19854 23714 19906 23726
rect 19854 23650 19906 23662
rect 26574 23714 26626 23726
rect 26574 23650 26626 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 23998 23266 24050 23278
rect 23998 23202 24050 23214
rect 25342 23266 25394 23278
rect 25342 23202 25394 23214
rect 25902 23266 25954 23278
rect 25902 23202 25954 23214
rect 22430 23154 22482 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 16482 23102 16494 23154
rect 16546 23102 16558 23154
rect 18946 23102 18958 23154
rect 19010 23102 19022 23154
rect 22430 23090 22482 23102
rect 24110 23154 24162 23166
rect 24110 23090 24162 23102
rect 25454 23154 25506 23166
rect 25454 23090 25506 23102
rect 25790 23154 25842 23166
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 25790 23090 25842 23102
rect 17502 23042 17554 23054
rect 21758 23042 21810 23054
rect 13682 22990 13694 23042
rect 13746 22990 13758 23042
rect 15810 22990 15822 23042
rect 15874 22990 15886 23042
rect 19618 22990 19630 23042
rect 19682 22990 19694 23042
rect 17502 22978 17554 22990
rect 21758 22978 21810 22990
rect 24334 23042 24386 23054
rect 24334 22978 24386 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 23550 22930 23602 22942
rect 23550 22866 23602 22878
rect 23774 22930 23826 22942
rect 23774 22866 23826 22878
rect 25342 22930 25394 22942
rect 25342 22866 25394 22878
rect 25902 22930 25954 22942
rect 25902 22866 25954 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 17726 22594 17778 22606
rect 17726 22530 17778 22542
rect 1934 22482 1986 22494
rect 13582 22482 13634 22494
rect 9986 22430 9998 22482
rect 10050 22430 10062 22482
rect 1934 22418 1986 22430
rect 13582 22418 13634 22430
rect 14590 22482 14642 22494
rect 19630 22482 19682 22494
rect 17378 22430 17390 22482
rect 17442 22430 17454 22482
rect 26226 22430 26238 22482
rect 26290 22430 26302 22482
rect 14590 22418 14642 22430
rect 19630 22418 19682 22430
rect 13918 22370 13970 22382
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 12898 22318 12910 22370
rect 12962 22318 12974 22370
rect 13918 22306 13970 22318
rect 14254 22370 14306 22382
rect 14254 22306 14306 22318
rect 15598 22370 15650 22382
rect 15598 22306 15650 22318
rect 16606 22370 16658 22382
rect 16606 22306 16658 22318
rect 16830 22370 16882 22382
rect 19854 22370 19906 22382
rect 26686 22370 26738 22382
rect 19282 22318 19294 22370
rect 19346 22318 19358 22370
rect 21410 22318 21422 22370
rect 21474 22318 21486 22370
rect 23314 22318 23326 22370
rect 23378 22318 23390 22370
rect 16830 22306 16882 22318
rect 19854 22306 19906 22318
rect 26686 22306 26738 22318
rect 14142 22258 14194 22270
rect 12114 22206 12126 22258
rect 12178 22206 12190 22258
rect 14142 22194 14194 22206
rect 15710 22258 15762 22270
rect 15710 22194 15762 22206
rect 16158 22258 16210 22270
rect 17054 22258 17106 22270
rect 16370 22206 16382 22258
rect 16434 22206 16446 22258
rect 16158 22194 16210 22206
rect 17054 22194 17106 22206
rect 17502 22258 17554 22270
rect 17502 22194 17554 22206
rect 19518 22258 19570 22270
rect 24098 22206 24110 22258
rect 24162 22206 24174 22258
rect 19518 22194 19570 22206
rect 14702 22146 14754 22158
rect 14702 22082 14754 22094
rect 15934 22146 15986 22158
rect 19742 22146 19794 22158
rect 16482 22094 16494 22146
rect 16546 22094 16558 22146
rect 21634 22094 21646 22146
rect 21698 22094 21710 22146
rect 15934 22082 15986 22094
rect 19742 22082 19794 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14702 21810 14754 21822
rect 14702 21746 14754 21758
rect 19630 21810 19682 21822
rect 22194 21758 22206 21810
rect 22258 21758 22270 21810
rect 19630 21746 19682 21758
rect 14814 21698 14866 21710
rect 19070 21698 19122 21710
rect 19854 21698 19906 21710
rect 18386 21646 18398 21698
rect 18450 21646 18462 21698
rect 19394 21646 19406 21698
rect 19458 21646 19470 21698
rect 14814 21634 14866 21646
rect 19070 21634 19122 21646
rect 19854 21634 19906 21646
rect 19966 21698 20018 21710
rect 24110 21698 24162 21710
rect 21522 21646 21534 21698
rect 21586 21646 21598 21698
rect 22082 21646 22094 21698
rect 22146 21646 22158 21698
rect 19966 21634 20018 21646
rect 24110 21634 24162 21646
rect 24446 21698 24498 21710
rect 24446 21634 24498 21646
rect 15038 21586 15090 21598
rect 15822 21586 15874 21598
rect 23886 21586 23938 21598
rect 15474 21534 15486 21586
rect 15538 21534 15550 21586
rect 18610 21534 18622 21586
rect 18674 21534 18686 21586
rect 21186 21534 21198 21586
rect 21250 21534 21262 21586
rect 15038 21522 15090 21534
rect 15822 21522 15874 21534
rect 23886 21522 23938 21534
rect 24222 21586 24274 21598
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 24222 21522 24274 21534
rect 18062 21474 18114 21486
rect 18062 21410 18114 21422
rect 15262 21362 15314 21374
rect 15262 21298 15314 21310
rect 23662 21362 23714 21374
rect 23662 21298 23714 21310
rect 40014 21362 40066 21374
rect 40014 21298 40066 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 25218 20862 25230 20914
rect 25282 20862 25294 20914
rect 21198 20802 21250 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 22642 20750 22654 20802
rect 22706 20750 22718 20802
rect 21198 20738 21250 20750
rect 21534 20690 21586 20702
rect 17042 20638 17054 20690
rect 17106 20638 17118 20690
rect 21534 20626 21586 20638
rect 21422 20578 21474 20590
rect 21422 20514 21474 20526
rect 21982 20578 22034 20590
rect 22194 20526 22206 20578
rect 22258 20575 22270 20578
rect 22530 20575 22542 20578
rect 22258 20529 22542 20575
rect 22258 20526 22270 20529
rect 22530 20526 22542 20529
rect 22594 20526 22606 20578
rect 21982 20514 22034 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 17838 20130 17890 20142
rect 15474 20078 15486 20130
rect 15538 20078 15550 20130
rect 16482 20078 16494 20130
rect 16546 20078 16558 20130
rect 17838 20066 17890 20078
rect 18510 20130 18562 20142
rect 22642 20078 22654 20130
rect 22706 20078 22718 20130
rect 18510 20066 18562 20078
rect 15822 20018 15874 20030
rect 15822 19954 15874 19966
rect 16158 20018 16210 20030
rect 16158 19954 16210 19966
rect 17614 20018 17666 20030
rect 17614 19954 17666 19966
rect 17950 20018 18002 20030
rect 17950 19954 18002 19966
rect 18286 20018 18338 20030
rect 29038 20018 29090 20030
rect 18946 19966 18958 20018
rect 19010 19966 19022 20018
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 18286 19954 18338 19966
rect 29038 19954 29090 19966
rect 29486 19906 29538 19918
rect 18610 19854 18622 19906
rect 18674 19854 18686 19906
rect 26450 19854 26462 19906
rect 26514 19854 26526 19906
rect 28578 19854 28590 19906
rect 28642 19854 28654 19906
rect 29486 19842 29538 19854
rect 28926 19794 28978 19806
rect 28926 19730 28978 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 15038 19458 15090 19470
rect 15038 19394 15090 19406
rect 15374 19458 15426 19470
rect 15374 19394 15426 19406
rect 15822 19458 15874 19470
rect 15822 19394 15874 19406
rect 17614 19458 17666 19470
rect 17614 19394 17666 19406
rect 1934 19346 1986 19358
rect 1934 19282 1986 19294
rect 15262 19346 15314 19358
rect 21422 19346 21474 19358
rect 27918 19346 27970 19358
rect 16594 19294 16606 19346
rect 16658 19294 16670 19346
rect 26898 19294 26910 19346
rect 26962 19294 26974 19346
rect 15262 19282 15314 19294
rect 21422 19282 21474 19294
rect 27918 19282 27970 19294
rect 14702 19234 14754 19246
rect 19294 19234 19346 19246
rect 4274 19182 4286 19234
rect 4338 19182 4350 19234
rect 18162 19182 18174 19234
rect 18226 19182 18238 19234
rect 18722 19182 18734 19234
rect 18786 19182 18798 19234
rect 14702 19170 14754 19182
rect 19294 19170 19346 19182
rect 19966 19234 20018 19246
rect 20750 19234 20802 19246
rect 20178 19182 20190 19234
rect 20242 19182 20254 19234
rect 19966 19170 20018 19182
rect 20750 19170 20802 19182
rect 22318 19234 22370 19246
rect 22318 19170 22370 19182
rect 22878 19234 22930 19246
rect 22878 19170 22930 19182
rect 23326 19234 23378 19246
rect 24098 19182 24110 19234
rect 24162 19182 24174 19234
rect 23326 19170 23378 19182
rect 14926 19122 14978 19134
rect 14926 19058 14978 19070
rect 15934 19122 15986 19134
rect 15934 19058 15986 19070
rect 16158 19122 16210 19134
rect 16158 19058 16210 19070
rect 16718 19122 16770 19134
rect 16718 19058 16770 19070
rect 16942 19122 16994 19134
rect 16942 19058 16994 19070
rect 18958 19122 19010 19134
rect 21310 19122 21362 19134
rect 19618 19070 19630 19122
rect 19682 19070 19694 19122
rect 18958 19058 19010 19070
rect 21310 19058 21362 19070
rect 21534 19122 21586 19134
rect 21534 19058 21586 19070
rect 22654 19122 22706 19134
rect 27358 19122 27410 19134
rect 24770 19070 24782 19122
rect 24834 19070 24846 19122
rect 22654 19058 22706 19070
rect 27358 19058 27410 19070
rect 27470 19122 27522 19134
rect 27470 19058 27522 19070
rect 14030 19010 14082 19022
rect 14030 18946 14082 18958
rect 14142 19010 14194 19022
rect 14142 18946 14194 18958
rect 14254 19010 14306 19022
rect 14254 18946 14306 18958
rect 17390 19010 17442 19022
rect 17390 18946 17442 18958
rect 17502 19010 17554 19022
rect 22542 19010 22594 19022
rect 27134 19010 27186 19022
rect 17938 18958 17950 19010
rect 18002 18958 18014 19010
rect 23650 18958 23662 19010
rect 23714 18958 23726 19010
rect 17502 18946 17554 18958
rect 22542 18946 22594 18958
rect 27134 18946 27186 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 17726 18674 17778 18686
rect 17726 18610 17778 18622
rect 21982 18674 22034 18686
rect 24222 18674 24274 18686
rect 22306 18622 22318 18674
rect 22370 18622 22382 18674
rect 21982 18610 22034 18622
rect 24222 18610 24274 18622
rect 24334 18674 24386 18686
rect 24334 18610 24386 18622
rect 24558 18674 24610 18686
rect 24558 18610 24610 18622
rect 26014 18674 26066 18686
rect 26014 18610 26066 18622
rect 26126 18674 26178 18686
rect 26126 18610 26178 18622
rect 26238 18674 26290 18686
rect 26238 18610 26290 18622
rect 14590 18562 14642 18574
rect 18062 18562 18114 18574
rect 16258 18510 16270 18562
rect 16322 18510 16334 18562
rect 14590 18498 14642 18510
rect 18062 18498 18114 18510
rect 19294 18562 19346 18574
rect 24110 18562 24162 18574
rect 19730 18510 19742 18562
rect 19794 18510 19806 18562
rect 20738 18510 20750 18562
rect 20802 18510 20814 18562
rect 22754 18510 22766 18562
rect 22818 18510 22830 18562
rect 23202 18510 23214 18562
rect 23266 18510 23278 18562
rect 19294 18498 19346 18510
rect 24110 18498 24162 18510
rect 27022 18562 27074 18574
rect 27022 18498 27074 18510
rect 14814 18450 14866 18462
rect 11106 18398 11118 18450
rect 11170 18398 11182 18450
rect 11778 18398 11790 18450
rect 11842 18398 11854 18450
rect 14814 18386 14866 18398
rect 15150 18450 15202 18462
rect 15150 18386 15202 18398
rect 15374 18450 15426 18462
rect 15374 18386 15426 18398
rect 15934 18450 15986 18462
rect 15934 18386 15986 18398
rect 17614 18450 17666 18462
rect 17614 18386 17666 18398
rect 18174 18450 18226 18462
rect 19070 18450 19122 18462
rect 26350 18450 26402 18462
rect 27246 18450 27298 18462
rect 18722 18398 18734 18450
rect 18786 18398 18798 18450
rect 19954 18398 19966 18450
rect 20018 18398 20030 18450
rect 20514 18398 20526 18450
rect 20578 18398 20590 18450
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 22306 18398 22318 18450
rect 22370 18398 22382 18450
rect 23426 18398 23438 18450
rect 23490 18398 23502 18450
rect 25778 18398 25790 18450
rect 25842 18398 25854 18450
rect 26786 18398 26798 18450
rect 26850 18398 26862 18450
rect 18174 18386 18226 18398
rect 19070 18386 19122 18398
rect 26350 18386 26402 18398
rect 27246 18386 27298 18398
rect 27358 18450 27410 18462
rect 27358 18386 27410 18398
rect 27134 18338 27186 18350
rect 13906 18286 13918 18338
rect 13970 18286 13982 18338
rect 27134 18274 27186 18286
rect 14702 18226 14754 18238
rect 14702 18162 14754 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 17950 17890 18002 17902
rect 13906 17838 13918 17890
rect 13970 17887 13982 17890
rect 14578 17887 14590 17890
rect 13970 17841 14590 17887
rect 13970 17838 13982 17841
rect 14578 17838 14590 17841
rect 14642 17838 14654 17890
rect 17950 17826 18002 17838
rect 23550 17890 23602 17902
rect 23550 17826 23602 17838
rect 25006 17890 25058 17902
rect 25006 17826 25058 17838
rect 21534 17778 21586 17790
rect 29262 17778 29314 17790
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 12114 17726 12126 17778
rect 12178 17726 12190 17778
rect 19842 17726 19854 17778
rect 19906 17726 19918 17778
rect 26450 17726 26462 17778
rect 26514 17726 26526 17778
rect 28578 17726 28590 17778
rect 28642 17726 28654 17778
rect 21534 17714 21586 17726
rect 29262 17714 29314 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 13582 17666 13634 17678
rect 12786 17614 12798 17666
rect 12850 17614 12862 17666
rect 13582 17602 13634 17614
rect 14142 17666 14194 17678
rect 14142 17602 14194 17614
rect 15150 17666 15202 17678
rect 15150 17602 15202 17614
rect 16158 17666 16210 17678
rect 16158 17602 16210 17614
rect 16494 17666 16546 17678
rect 16494 17602 16546 17614
rect 16718 17666 16770 17678
rect 18062 17666 18114 17678
rect 17602 17614 17614 17666
rect 17666 17614 17678 17666
rect 19170 17614 19182 17666
rect 19234 17614 19246 17666
rect 20290 17614 20302 17666
rect 20354 17614 20366 17666
rect 24658 17614 24670 17666
rect 24722 17614 24734 17666
rect 25666 17614 25678 17666
rect 25730 17614 25742 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 16718 17602 16770 17614
rect 18062 17602 18114 17614
rect 15486 17554 15538 17566
rect 14802 17502 14814 17554
rect 14866 17502 14878 17554
rect 15486 17490 15538 17502
rect 15822 17554 15874 17566
rect 15822 17490 15874 17502
rect 18398 17554 18450 17566
rect 21422 17554 21474 17566
rect 20066 17502 20078 17554
rect 20130 17502 20142 17554
rect 18398 17490 18450 17502
rect 21422 17490 21474 17502
rect 21646 17554 21698 17566
rect 21646 17490 21698 17502
rect 23438 17554 23490 17566
rect 23438 17490 23490 17502
rect 23550 17554 23602 17566
rect 23550 17490 23602 17502
rect 24110 17554 24162 17566
rect 24110 17490 24162 17502
rect 24446 17554 24498 17566
rect 24446 17490 24498 17502
rect 24894 17554 24946 17566
rect 24894 17490 24946 17502
rect 16494 17442 16546 17454
rect 17938 17390 17950 17442
rect 18002 17390 18014 17442
rect 16494 17378 16546 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 17614 17106 17666 17118
rect 17614 17042 17666 17054
rect 20078 17106 20130 17118
rect 20078 17042 20130 17054
rect 20526 17106 20578 17118
rect 27694 17106 27746 17118
rect 20850 17054 20862 17106
rect 20914 17054 20926 17106
rect 21186 17054 21198 17106
rect 21250 17054 21262 17106
rect 20526 17042 20578 17054
rect 27694 17042 27746 17054
rect 13918 16994 13970 17006
rect 13918 16930 13970 16942
rect 19966 16994 20018 17006
rect 19966 16930 20018 16942
rect 20302 16994 20354 17006
rect 26686 16994 26738 17006
rect 22306 16942 22318 16994
rect 22370 16942 22382 16994
rect 20302 16930 20354 16942
rect 26686 16930 26738 16942
rect 27246 16994 27298 17006
rect 27246 16930 27298 16942
rect 27358 16994 27410 17006
rect 27358 16930 27410 16942
rect 27806 16994 27858 17006
rect 27806 16930 27858 16942
rect 14030 16882 14082 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 14030 16818 14082 16830
rect 14254 16882 14306 16894
rect 26462 16882 26514 16894
rect 14690 16830 14702 16882
rect 14754 16830 14766 16882
rect 21410 16830 21422 16882
rect 21474 16830 21486 16882
rect 22530 16830 22542 16882
rect 22594 16830 22606 16882
rect 14254 16818 14306 16830
rect 26462 16818 26514 16830
rect 26798 16882 26850 16894
rect 26798 16818 26850 16830
rect 27022 16882 27074 16894
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 27022 16818 27074 16830
rect 14366 16770 14418 16782
rect 14366 16706 14418 16718
rect 17390 16770 17442 16782
rect 17390 16706 17442 16718
rect 17502 16770 17554 16782
rect 17502 16706 17554 16718
rect 40014 16770 40066 16782
rect 40014 16706 40066 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 14254 16322 14306 16334
rect 14254 16258 14306 16270
rect 15598 16322 15650 16334
rect 15598 16258 15650 16270
rect 29262 16210 29314 16222
rect 2034 16158 2046 16210
rect 2098 16158 2110 16210
rect 15250 16158 15262 16210
rect 15314 16158 15326 16210
rect 21858 16158 21870 16210
rect 21922 16158 21934 16210
rect 26450 16158 26462 16210
rect 26514 16158 26526 16210
rect 28578 16158 28590 16210
rect 28642 16158 28654 16210
rect 29262 16146 29314 16158
rect 18286 16098 18338 16110
rect 4050 16046 4062 16098
rect 4114 16046 4126 16098
rect 13682 16046 13694 16098
rect 13746 16046 13758 16098
rect 18286 16034 18338 16046
rect 18622 16098 18674 16110
rect 18622 16034 18674 16046
rect 18734 16098 18786 16110
rect 19518 16098 19570 16110
rect 19966 16098 20018 16110
rect 22318 16098 22370 16110
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 19730 16046 19742 16098
rect 19794 16046 19806 16098
rect 20514 16046 20526 16098
rect 20578 16046 20590 16098
rect 24210 16046 24222 16098
rect 24274 16046 24286 16098
rect 25666 16046 25678 16098
rect 25730 16046 25742 16098
rect 18734 16034 18786 16046
rect 19518 16034 19570 16046
rect 19966 16034 20018 16046
rect 22318 16034 22370 16046
rect 14142 15986 14194 15998
rect 14142 15922 14194 15934
rect 15374 15986 15426 15998
rect 24446 15986 24498 15998
rect 20290 15934 20302 15986
rect 20354 15934 20366 15986
rect 22978 15934 22990 15986
rect 23042 15934 23054 15986
rect 15374 15922 15426 15934
rect 24446 15922 24498 15934
rect 18398 15874 18450 15886
rect 13458 15822 13470 15874
rect 13522 15822 13534 15874
rect 18398 15810 18450 15822
rect 19182 15874 19234 15886
rect 19182 15810 19234 15822
rect 22654 15874 22706 15886
rect 22654 15810 22706 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 20414 15538 20466 15550
rect 20414 15474 20466 15486
rect 22430 15538 22482 15550
rect 22430 15474 22482 15486
rect 19518 15426 19570 15438
rect 12786 15374 12798 15426
rect 12850 15374 12862 15426
rect 14690 15374 14702 15426
rect 14754 15374 14766 15426
rect 19518 15362 19570 15374
rect 24222 15426 24274 15438
rect 24222 15362 24274 15374
rect 17502 15314 17554 15326
rect 4274 15262 4286 15314
rect 4338 15262 4350 15314
rect 13570 15262 13582 15314
rect 13634 15262 13646 15314
rect 13906 15262 13918 15314
rect 13970 15262 13982 15314
rect 17502 15250 17554 15262
rect 19630 15314 19682 15326
rect 20190 15314 20242 15326
rect 19954 15262 19966 15314
rect 20018 15262 20030 15314
rect 19630 15250 19682 15262
rect 20190 15250 20242 15262
rect 20526 15314 20578 15326
rect 23326 15314 23378 15326
rect 22194 15262 22206 15314
rect 22258 15262 22270 15314
rect 23538 15262 23550 15314
rect 23602 15262 23614 15314
rect 20526 15250 20578 15262
rect 23326 15250 23378 15262
rect 10658 15150 10670 15202
rect 10722 15150 10734 15202
rect 16818 15150 16830 15202
rect 16882 15150 16894 15202
rect 20066 15150 20078 15202
rect 20130 15150 20142 15202
rect 1934 15090 1986 15102
rect 1934 15026 1986 15038
rect 22542 15090 22594 15102
rect 22542 15026 22594 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 14254 14642 14306 14654
rect 26910 14642 26962 14654
rect 23090 14590 23102 14642
rect 23154 14590 23166 14642
rect 23538 14590 23550 14642
rect 23602 14590 23614 14642
rect 14254 14578 14306 14590
rect 26910 14578 26962 14590
rect 18286 14530 18338 14542
rect 13682 14478 13694 14530
rect 13746 14478 13758 14530
rect 18286 14466 18338 14478
rect 21534 14530 21586 14542
rect 21534 14466 21586 14478
rect 21982 14530 22034 14542
rect 26338 14478 26350 14530
rect 26402 14478 26414 14530
rect 21982 14466 22034 14478
rect 17838 14418 17890 14430
rect 22306 14366 22318 14418
rect 22370 14366 22382 14418
rect 25666 14366 25678 14418
rect 25730 14366 25742 14418
rect 17838 14354 17890 14366
rect 18062 14306 18114 14318
rect 13458 14254 13470 14306
rect 13522 14254 13534 14306
rect 18062 14242 18114 14254
rect 18174 14306 18226 14318
rect 18174 14242 18226 14254
rect 21646 14306 21698 14318
rect 21646 14242 21698 14254
rect 22654 14306 22706 14318
rect 22654 14242 22706 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 17614 13970 17666 13982
rect 17614 13906 17666 13918
rect 18722 13806 18734 13858
rect 18786 13806 18798 13858
rect 23314 13806 23326 13858
rect 23378 13806 23390 13858
rect 24558 13746 24610 13758
rect 17938 13694 17950 13746
rect 18002 13694 18014 13746
rect 24098 13694 24110 13746
rect 24162 13694 24174 13746
rect 24558 13682 24610 13694
rect 17502 13634 17554 13646
rect 20850 13582 20862 13634
rect 20914 13582 20926 13634
rect 21186 13582 21198 13634
rect 21250 13582 21262 13634
rect 17502 13570 17554 13582
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 19182 13074 19234 13086
rect 15810 13022 15822 13074
rect 15874 13022 15886 13074
rect 17938 13022 17950 13074
rect 18002 13022 18014 13074
rect 19182 13010 19234 13022
rect 18610 12910 18622 12962
rect 18674 12910 18686 12962
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 15374 38222 15426 38274
rect 19182 38222 19234 38274
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 15934 37998 15986 38050
rect 19742 37998 19794 38050
rect 21422 37998 21474 38050
rect 25006 37998 25058 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 22766 37438 22818 37490
rect 26238 37438 26290 37490
rect 21198 37214 21250 37266
rect 21870 37214 21922 37266
rect 25566 37214 25618 37266
rect 20078 37102 20130 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 18062 36654 18114 36706
rect 22318 36654 22370 36706
rect 26126 36654 26178 36706
rect 17166 36430 17218 36482
rect 21758 36430 21810 36482
rect 25230 36430 25282 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 14478 28366 14530 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 14814 28030 14866 28082
rect 14142 27806 14194 27858
rect 15038 27806 15090 27858
rect 15374 27806 15426 27858
rect 15598 27806 15650 27858
rect 16046 27806 16098 27858
rect 18958 27806 19010 27858
rect 22318 27806 22370 27858
rect 11230 27694 11282 27746
rect 13358 27694 13410 27746
rect 17502 27694 17554 27746
rect 19630 27694 19682 27746
rect 21758 27694 21810 27746
rect 15150 27582 15202 27634
rect 15934 27582 15986 27634
rect 16046 27582 16098 27634
rect 16494 27582 16546 27634
rect 16718 27582 16770 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1934 27134 1986 27186
rect 15038 27134 15090 27186
rect 17166 27134 17218 27186
rect 20526 27134 20578 27186
rect 25006 27134 25058 27186
rect 4286 27022 4338 27074
rect 14254 27022 14306 27074
rect 17614 27022 17666 27074
rect 22206 27022 22258 27074
rect 25678 27022 25730 27074
rect 18398 26910 18450 26962
rect 21310 26910 21362 26962
rect 21422 26910 21474 26962
rect 21646 26910 21698 26962
rect 22878 26910 22930 26962
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 16158 26462 16210 26514
rect 16270 26462 16322 26514
rect 18734 26462 18786 26514
rect 19742 26462 19794 26514
rect 20750 26462 20802 26514
rect 22318 26462 22370 26514
rect 23662 26462 23714 26514
rect 24334 26462 24386 26514
rect 24670 26462 24722 26514
rect 25230 26462 25282 26514
rect 25566 26462 25618 26514
rect 13806 26350 13858 26402
rect 19518 26350 19570 26402
rect 19966 26350 20018 26402
rect 21310 26350 21362 26402
rect 21646 26350 21698 26402
rect 22430 26350 22482 26402
rect 13134 26238 13186 26290
rect 16494 26238 16546 26290
rect 16830 26238 16882 26290
rect 18510 26238 18562 26290
rect 18846 26238 18898 26290
rect 19182 26238 19234 26290
rect 20414 26238 20466 26290
rect 20750 26238 20802 26290
rect 21086 26238 21138 26290
rect 22206 26238 22258 26290
rect 22878 26238 22930 26290
rect 23438 26238 23490 26290
rect 23774 26238 23826 26290
rect 15934 26126 15986 26178
rect 17502 26126 17554 26178
rect 19630 26126 19682 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 14814 25678 14866 25730
rect 15710 25678 15762 25730
rect 15822 25566 15874 25618
rect 14142 25342 14194 25394
rect 14254 25342 14306 25394
rect 14478 25342 14530 25394
rect 14702 25342 14754 25394
rect 15150 25342 15202 25394
rect 19854 25342 19906 25394
rect 14926 25230 14978 25282
rect 16270 25230 16322 25282
rect 20190 25230 20242 25282
rect 20638 25230 20690 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 17614 24894 17666 24946
rect 20750 24894 20802 24946
rect 21086 24894 21138 24946
rect 13918 24670 13970 24722
rect 14366 24670 14418 24722
rect 17838 24670 17890 24722
rect 11006 24558 11058 24610
rect 13134 24558 13186 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 1934 23998 1986 24050
rect 15934 23998 15986 24050
rect 19518 23998 19570 24050
rect 26126 23998 26178 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 15486 23886 15538 23938
rect 16158 23886 16210 23938
rect 16718 23886 16770 23938
rect 21422 23886 21474 23938
rect 23214 23886 23266 23938
rect 37886 23886 37938 23938
rect 14366 23774 14418 23826
rect 14478 23774 14530 23826
rect 15710 23774 15762 23826
rect 17278 23774 17330 23826
rect 19406 23774 19458 23826
rect 21646 23774 21698 23826
rect 23998 23774 24050 23826
rect 14142 23662 14194 23714
rect 15598 23662 15650 23714
rect 16494 23662 16546 23714
rect 19630 23662 19682 23714
rect 19854 23662 19906 23714
rect 26574 23662 26626 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 23998 23214 24050 23266
rect 25342 23214 25394 23266
rect 25902 23214 25954 23266
rect 4286 23102 4338 23154
rect 16494 23102 16546 23154
rect 18958 23102 19010 23154
rect 22430 23102 22482 23154
rect 24110 23102 24162 23154
rect 25454 23102 25506 23154
rect 25790 23102 25842 23154
rect 37662 23102 37714 23154
rect 13694 22990 13746 23042
rect 15822 22990 15874 23042
rect 17502 22990 17554 23042
rect 19630 22990 19682 23042
rect 21758 22990 21810 23042
rect 24334 22990 24386 23042
rect 1934 22878 1986 22930
rect 23550 22878 23602 22930
rect 23774 22878 23826 22930
rect 25342 22878 25394 22930
rect 25902 22878 25954 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 17726 22542 17778 22594
rect 1934 22430 1986 22482
rect 9998 22430 10050 22482
rect 13582 22430 13634 22482
rect 14590 22430 14642 22482
rect 17390 22430 17442 22482
rect 19630 22430 19682 22482
rect 26238 22430 26290 22482
rect 4286 22318 4338 22370
rect 12910 22318 12962 22370
rect 13918 22318 13970 22370
rect 14254 22318 14306 22370
rect 15598 22318 15650 22370
rect 16606 22318 16658 22370
rect 16830 22318 16882 22370
rect 19294 22318 19346 22370
rect 19854 22318 19906 22370
rect 21422 22318 21474 22370
rect 23326 22318 23378 22370
rect 26686 22318 26738 22370
rect 12126 22206 12178 22258
rect 14142 22206 14194 22258
rect 15710 22206 15762 22258
rect 16158 22206 16210 22258
rect 16382 22206 16434 22258
rect 17054 22206 17106 22258
rect 17502 22206 17554 22258
rect 19518 22206 19570 22258
rect 24110 22206 24162 22258
rect 14702 22094 14754 22146
rect 15934 22094 15986 22146
rect 16494 22094 16546 22146
rect 19742 22094 19794 22146
rect 21646 22094 21698 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14702 21758 14754 21810
rect 19630 21758 19682 21810
rect 22206 21758 22258 21810
rect 14814 21646 14866 21698
rect 18398 21646 18450 21698
rect 19070 21646 19122 21698
rect 19406 21646 19458 21698
rect 19854 21646 19906 21698
rect 19966 21646 20018 21698
rect 21534 21646 21586 21698
rect 22094 21646 22146 21698
rect 24110 21646 24162 21698
rect 24446 21646 24498 21698
rect 15038 21534 15090 21586
rect 15486 21534 15538 21586
rect 15822 21534 15874 21586
rect 18622 21534 18674 21586
rect 21198 21534 21250 21586
rect 23886 21534 23938 21586
rect 24222 21534 24274 21586
rect 37886 21534 37938 21586
rect 18062 21422 18114 21474
rect 15262 21310 15314 21362
rect 23662 21310 23714 21362
rect 40014 21310 40066 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 25230 20862 25282 20914
rect 20078 20750 20130 20802
rect 21198 20750 21250 20802
rect 22654 20750 22706 20802
rect 17054 20638 17106 20690
rect 21534 20638 21586 20690
rect 21422 20526 21474 20578
rect 21982 20526 22034 20578
rect 22206 20526 22258 20578
rect 22542 20526 22594 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 15486 20078 15538 20130
rect 16494 20078 16546 20130
rect 17838 20078 17890 20130
rect 18510 20078 18562 20130
rect 22654 20078 22706 20130
rect 15822 19966 15874 20018
rect 16158 19966 16210 20018
rect 17614 19966 17666 20018
rect 17950 19966 18002 20018
rect 18286 19966 18338 20018
rect 18958 19966 19010 20018
rect 25678 19966 25730 20018
rect 29038 19966 29090 20018
rect 37662 19966 37714 20018
rect 18622 19854 18674 19906
rect 26462 19854 26514 19906
rect 28590 19854 28642 19906
rect 29486 19854 29538 19906
rect 28926 19742 28978 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15038 19406 15090 19458
rect 15374 19406 15426 19458
rect 15822 19406 15874 19458
rect 17614 19406 17666 19458
rect 1934 19294 1986 19346
rect 15262 19294 15314 19346
rect 16606 19294 16658 19346
rect 21422 19294 21474 19346
rect 26910 19294 26962 19346
rect 27918 19294 27970 19346
rect 4286 19182 4338 19234
rect 14702 19182 14754 19234
rect 18174 19182 18226 19234
rect 18734 19182 18786 19234
rect 19294 19182 19346 19234
rect 19966 19182 20018 19234
rect 20190 19182 20242 19234
rect 20750 19182 20802 19234
rect 22318 19182 22370 19234
rect 22878 19182 22930 19234
rect 23326 19182 23378 19234
rect 24110 19182 24162 19234
rect 14926 19070 14978 19122
rect 15934 19070 15986 19122
rect 16158 19070 16210 19122
rect 16718 19070 16770 19122
rect 16942 19070 16994 19122
rect 18958 19070 19010 19122
rect 19630 19070 19682 19122
rect 21310 19070 21362 19122
rect 21534 19070 21586 19122
rect 22654 19070 22706 19122
rect 24782 19070 24834 19122
rect 27358 19070 27410 19122
rect 27470 19070 27522 19122
rect 14030 18958 14082 19010
rect 14142 18958 14194 19010
rect 14254 18958 14306 19010
rect 17390 18958 17442 19010
rect 17502 18958 17554 19010
rect 17950 18958 18002 19010
rect 22542 18958 22594 19010
rect 23662 18958 23714 19010
rect 27134 18958 27186 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 17726 18622 17778 18674
rect 21982 18622 22034 18674
rect 22318 18622 22370 18674
rect 24222 18622 24274 18674
rect 24334 18622 24386 18674
rect 24558 18622 24610 18674
rect 26014 18622 26066 18674
rect 26126 18622 26178 18674
rect 26238 18622 26290 18674
rect 14590 18510 14642 18562
rect 16270 18510 16322 18562
rect 18062 18510 18114 18562
rect 19294 18510 19346 18562
rect 19742 18510 19794 18562
rect 20750 18510 20802 18562
rect 22766 18510 22818 18562
rect 23214 18510 23266 18562
rect 24110 18510 24162 18562
rect 27022 18510 27074 18562
rect 11118 18398 11170 18450
rect 11790 18398 11842 18450
rect 14814 18398 14866 18450
rect 15150 18398 15202 18450
rect 15374 18398 15426 18450
rect 15934 18398 15986 18450
rect 17614 18398 17666 18450
rect 18174 18398 18226 18450
rect 18734 18398 18786 18450
rect 19070 18398 19122 18450
rect 19966 18398 20018 18450
rect 20526 18398 20578 18450
rect 21422 18398 21474 18450
rect 22318 18398 22370 18450
rect 23438 18398 23490 18450
rect 25790 18398 25842 18450
rect 26350 18398 26402 18450
rect 26798 18398 26850 18450
rect 27246 18398 27298 18450
rect 27358 18398 27410 18450
rect 13918 18286 13970 18338
rect 27134 18286 27186 18338
rect 14702 18174 14754 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 13918 17838 13970 17890
rect 14590 17838 14642 17890
rect 17950 17838 18002 17890
rect 23550 17838 23602 17890
rect 25006 17838 25058 17890
rect 9998 17726 10050 17778
rect 12126 17726 12178 17778
rect 19854 17726 19906 17778
rect 21534 17726 21586 17778
rect 26462 17726 26514 17778
rect 28590 17726 28642 17778
rect 29262 17726 29314 17778
rect 40014 17726 40066 17778
rect 12798 17614 12850 17666
rect 13582 17614 13634 17666
rect 14142 17614 14194 17666
rect 15150 17614 15202 17666
rect 16158 17614 16210 17666
rect 16494 17614 16546 17666
rect 16718 17614 16770 17666
rect 17614 17614 17666 17666
rect 18062 17614 18114 17666
rect 19182 17614 19234 17666
rect 20302 17614 20354 17666
rect 24670 17614 24722 17666
rect 25678 17614 25730 17666
rect 37662 17614 37714 17666
rect 14814 17502 14866 17554
rect 15486 17502 15538 17554
rect 15822 17502 15874 17554
rect 18398 17502 18450 17554
rect 20078 17502 20130 17554
rect 21422 17502 21474 17554
rect 21646 17502 21698 17554
rect 23438 17502 23490 17554
rect 23550 17502 23602 17554
rect 24110 17502 24162 17554
rect 24446 17502 24498 17554
rect 24894 17502 24946 17554
rect 16494 17390 16546 17442
rect 17950 17390 18002 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17614 17054 17666 17106
rect 20078 17054 20130 17106
rect 20526 17054 20578 17106
rect 20862 17054 20914 17106
rect 21198 17054 21250 17106
rect 27694 17054 27746 17106
rect 13918 16942 13970 16994
rect 19966 16942 20018 16994
rect 20302 16942 20354 16994
rect 22318 16942 22370 16994
rect 26686 16942 26738 16994
rect 27246 16942 27298 16994
rect 27358 16942 27410 16994
rect 27806 16942 27858 16994
rect 4286 16830 4338 16882
rect 14030 16830 14082 16882
rect 14254 16830 14306 16882
rect 14702 16830 14754 16882
rect 21422 16830 21474 16882
rect 22542 16830 22594 16882
rect 26462 16830 26514 16882
rect 26798 16830 26850 16882
rect 27022 16830 27074 16882
rect 37662 16830 37714 16882
rect 14366 16718 14418 16770
rect 17390 16718 17442 16770
rect 17502 16718 17554 16770
rect 40014 16718 40066 16770
rect 1934 16606 1986 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 14254 16270 14306 16322
rect 15598 16270 15650 16322
rect 2046 16158 2098 16210
rect 15262 16158 15314 16210
rect 21870 16158 21922 16210
rect 26462 16158 26514 16210
rect 28590 16158 28642 16210
rect 29262 16158 29314 16210
rect 4062 16046 4114 16098
rect 13694 16046 13746 16098
rect 18286 16046 18338 16098
rect 18622 16046 18674 16098
rect 18734 16046 18786 16098
rect 19182 16046 19234 16098
rect 19518 16046 19570 16098
rect 19742 16046 19794 16098
rect 19966 16046 20018 16098
rect 20526 16046 20578 16098
rect 22318 16046 22370 16098
rect 24222 16046 24274 16098
rect 25678 16046 25730 16098
rect 14142 15934 14194 15986
rect 15374 15934 15426 15986
rect 20302 15934 20354 15986
rect 22990 15934 23042 15986
rect 24446 15934 24498 15986
rect 13470 15822 13522 15874
rect 18398 15822 18450 15874
rect 19182 15822 19234 15874
rect 22654 15822 22706 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 20414 15486 20466 15538
rect 22430 15486 22482 15538
rect 12798 15374 12850 15426
rect 14702 15374 14754 15426
rect 19518 15374 19570 15426
rect 24222 15374 24274 15426
rect 4286 15262 4338 15314
rect 13582 15262 13634 15314
rect 13918 15262 13970 15314
rect 17502 15262 17554 15314
rect 19630 15262 19682 15314
rect 19966 15262 20018 15314
rect 20190 15262 20242 15314
rect 20526 15262 20578 15314
rect 22206 15262 22258 15314
rect 23326 15262 23378 15314
rect 23550 15262 23602 15314
rect 10670 15150 10722 15202
rect 16830 15150 16882 15202
rect 20078 15150 20130 15202
rect 1934 15038 1986 15090
rect 22542 15038 22594 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 14254 14590 14306 14642
rect 23102 14590 23154 14642
rect 23550 14590 23602 14642
rect 26910 14590 26962 14642
rect 13694 14478 13746 14530
rect 18286 14478 18338 14530
rect 21534 14478 21586 14530
rect 21982 14478 22034 14530
rect 26350 14478 26402 14530
rect 17838 14366 17890 14418
rect 22318 14366 22370 14418
rect 25678 14366 25730 14418
rect 13470 14254 13522 14306
rect 18062 14254 18114 14306
rect 18174 14254 18226 14306
rect 21646 14254 21698 14306
rect 22654 14254 22706 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 16830 13918 16882 13970
rect 17614 13918 17666 13970
rect 18734 13806 18786 13858
rect 23326 13806 23378 13858
rect 17950 13694 18002 13746
rect 24110 13694 24162 13746
rect 24558 13694 24610 13746
rect 17502 13582 17554 13634
rect 20862 13582 20914 13634
rect 21198 13582 21250 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 15822 13022 15874 13074
rect 17950 13022 18002 13074
rect 19182 13022 19234 13074
rect 18622 12910 18674 12962
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18622 3614 18674 3666
rect 22094 3614 22146 3666
rect 17614 3502 17666 3554
rect 21086 3502 21138 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16128 41200 16240 42000
rect 16800 41200 16912 42000
rect 19488 41200 19600 42000
rect 20160 41200 20272 42000
rect 20832 41200 20944 42000
rect 21504 41200 21616 42000
rect 22176 41200 22288 42000
rect 23520 41200 23632 42000
rect 24192 41200 24304 42000
rect 24864 41200 24976 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 15372 38276 15428 38286
rect 15372 38182 15428 38220
rect 16156 38276 16212 41200
rect 16156 38210 16212 38220
rect 15932 38050 15988 38062
rect 15932 37998 15934 38050
rect 15986 37998 15988 38050
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 15932 31948 15988 37998
rect 16828 36708 16884 41200
rect 19180 38276 19236 38286
rect 19516 38276 19572 41200
rect 19180 38274 19572 38276
rect 19180 38222 19182 38274
rect 19234 38222 19572 38274
rect 19180 38220 19572 38222
rect 19180 38210 19236 38220
rect 19740 38052 19796 38062
rect 19516 38050 19796 38052
rect 19516 37998 19742 38050
rect 19794 37998 19796 38050
rect 19516 37996 19796 37998
rect 16828 36642 16884 36652
rect 18060 36708 18116 36718
rect 18060 36614 18116 36652
rect 15820 31892 15988 31948
rect 17164 36482 17220 36494
rect 17164 36430 17166 36482
rect 17218 36430 17220 36482
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 14476 28418 14532 28430
rect 14476 28366 14478 28418
rect 14530 28366 14532 28418
rect 13804 28084 13860 28094
rect 11228 27746 11284 27758
rect 11228 27694 11230 27746
rect 11282 27694 11284 27746
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 4284 27076 4340 27086
rect 4284 26982 4340 27020
rect 11228 27076 11284 27694
rect 11228 27010 11284 27020
rect 13356 27746 13412 27758
rect 13356 27694 13358 27746
rect 13410 27694 13412 27746
rect 1932 26226 1988 26236
rect 4172 26964 4228 26974
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 1932 22484 1988 22494
rect 1932 22390 1988 22428
rect 4172 21476 4228 26908
rect 13132 26852 13188 26862
rect 13132 26290 13188 26796
rect 13132 26238 13134 26290
rect 13186 26238 13188 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13132 25284 13188 26238
rect 13356 25732 13412 27694
rect 13804 26402 13860 28028
rect 14140 27860 14196 27870
rect 14476 27860 14532 28366
rect 14812 28084 14868 28094
rect 14812 27990 14868 28028
rect 14140 27858 14532 27860
rect 14140 27806 14142 27858
rect 14194 27806 14532 27858
rect 14140 27804 14532 27806
rect 15036 27860 15092 27898
rect 14140 27794 14196 27804
rect 14140 27076 14196 27086
rect 14140 26740 14196 27020
rect 14252 27074 14308 27804
rect 15036 27794 15092 27804
rect 15372 27860 15428 27870
rect 15372 27858 15540 27860
rect 15372 27806 15374 27858
rect 15426 27806 15540 27858
rect 15372 27804 15540 27806
rect 15372 27794 15428 27804
rect 15036 27636 15092 27646
rect 15036 27186 15092 27580
rect 15036 27134 15038 27186
rect 15090 27134 15092 27186
rect 15036 27122 15092 27134
rect 15148 27634 15204 27646
rect 15148 27582 15150 27634
rect 15202 27582 15204 27634
rect 14252 27022 14254 27074
rect 14306 27022 14308 27074
rect 14252 26964 14308 27022
rect 14252 26898 14308 26908
rect 14140 26684 14308 26740
rect 13804 26350 13806 26402
rect 13858 26350 13860 26402
rect 13804 26338 13860 26350
rect 13356 25666 13412 25676
rect 14140 25396 14196 25406
rect 14140 25302 14196 25340
rect 14252 25394 14308 26684
rect 14812 25732 14868 25742
rect 14812 25638 14868 25676
rect 15148 25732 15204 27582
rect 15484 25732 15540 27804
rect 15596 27858 15652 27870
rect 15596 27806 15598 27858
rect 15650 27806 15652 27858
rect 15596 26852 15652 27806
rect 15596 26786 15652 26796
rect 15820 26180 15876 31892
rect 16044 27860 16100 27898
rect 16100 27804 16212 27860
rect 16044 27794 16100 27804
rect 15932 27634 15988 27646
rect 15932 27582 15934 27634
rect 15986 27582 15988 27634
rect 15932 26516 15988 27582
rect 16044 27636 16100 27646
rect 16044 27542 16100 27580
rect 16156 26740 16212 27804
rect 16492 27636 16548 27646
rect 16492 27634 16660 27636
rect 16492 27582 16494 27634
rect 16546 27582 16660 27634
rect 16492 27580 16660 27582
rect 16492 27570 16548 27580
rect 16156 26674 16212 26684
rect 16268 27188 16324 27198
rect 16156 26516 16212 26526
rect 15932 26514 16212 26516
rect 15932 26462 16158 26514
rect 16210 26462 16212 26514
rect 15932 26460 16212 26462
rect 16156 26450 16212 26460
rect 16268 26514 16324 27132
rect 16268 26462 16270 26514
rect 16322 26462 16324 26514
rect 16268 26450 16324 26462
rect 16604 26852 16660 27580
rect 16492 26290 16548 26302
rect 16492 26238 16494 26290
rect 16546 26238 16548 26290
rect 15932 26180 15988 26190
rect 15820 26178 15988 26180
rect 15820 26126 15934 26178
rect 15986 26126 15988 26178
rect 15820 26124 15988 26126
rect 15708 25732 15764 25742
rect 15484 25730 15764 25732
rect 15484 25678 15710 25730
rect 15762 25678 15764 25730
rect 15484 25676 15764 25678
rect 15148 25666 15204 25676
rect 15708 25666 15764 25676
rect 15372 25620 15428 25630
rect 15428 25564 15540 25620
rect 15372 25554 15428 25564
rect 15148 25508 15204 25518
rect 14252 25342 14254 25394
rect 14306 25342 14308 25394
rect 14252 25330 14308 25342
rect 14476 25396 14532 25406
rect 14700 25396 14756 25406
rect 14476 25394 14756 25396
rect 14476 25342 14478 25394
rect 14530 25342 14702 25394
rect 14754 25342 14756 25394
rect 14476 25340 14756 25342
rect 14476 25330 14532 25340
rect 14700 25330 14756 25340
rect 14812 25396 14868 25406
rect 13132 25218 13188 25228
rect 14364 25284 14420 25294
rect 13916 24724 13972 24734
rect 14364 24724 14420 25228
rect 13916 24722 14420 24724
rect 13916 24670 13918 24722
rect 13970 24670 14366 24722
rect 14418 24670 14420 24722
rect 13916 24668 14420 24670
rect 11004 24610 11060 24622
rect 11004 24558 11006 24610
rect 11058 24558 11060 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 11004 23828 11060 24558
rect 11004 23762 11060 23772
rect 13132 24610 13188 24622
rect 13132 24558 13134 24610
rect 13186 24558 13188 24610
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 13132 22596 13188 24558
rect 13692 23156 13748 23166
rect 13132 22530 13188 22540
rect 13580 23044 13636 23054
rect 9996 22484 10052 22494
rect 9996 22390 10052 22428
rect 13580 22482 13636 22988
rect 13692 23042 13748 23100
rect 13692 22990 13694 23042
rect 13746 22990 13748 23042
rect 13692 22978 13748 22990
rect 13916 23044 13972 24668
rect 14364 24658 14420 24668
rect 14364 23828 14420 23838
rect 14364 23734 14420 23772
rect 14476 23826 14532 23838
rect 14476 23774 14478 23826
rect 14530 23774 14532 23826
rect 13916 22978 13972 22988
rect 14140 23714 14196 23726
rect 14140 23662 14142 23714
rect 14194 23662 14196 23714
rect 13580 22430 13582 22482
rect 13634 22430 13636 22482
rect 4284 22372 4340 22382
rect 4284 22278 4340 22316
rect 12908 22372 12964 22382
rect 12908 22278 12964 22316
rect 13580 22372 13636 22430
rect 13580 22306 13636 22316
rect 13916 22596 13972 22606
rect 13916 22370 13972 22540
rect 13916 22318 13918 22370
rect 13970 22318 13972 22370
rect 13916 22306 13972 22318
rect 12124 22258 12180 22270
rect 12124 22206 12126 22258
rect 12178 22206 12180 22258
rect 12124 21812 12180 22206
rect 14140 22258 14196 23662
rect 14252 23716 14308 23726
rect 14252 22370 14308 23660
rect 14252 22318 14254 22370
rect 14306 22318 14308 22370
rect 14252 22306 14308 22318
rect 14476 22372 14532 23774
rect 14812 23828 14868 25340
rect 15148 25394 15204 25452
rect 15148 25342 15150 25394
rect 15202 25342 15204 25394
rect 15148 25330 15204 25342
rect 14924 25282 14980 25294
rect 14924 25230 14926 25282
rect 14978 25230 14980 25282
rect 14924 24052 14980 25230
rect 14924 23986 14980 23996
rect 15484 23940 15540 25564
rect 15820 25618 15876 26124
rect 15932 26114 15988 26124
rect 15820 25566 15822 25618
rect 15874 25566 15876 25618
rect 15820 25554 15876 25566
rect 16492 25396 16548 26238
rect 16604 26180 16660 26796
rect 16716 27634 16772 27646
rect 16716 27582 16718 27634
rect 16770 27582 16772 27634
rect 16716 26516 16772 27582
rect 17164 27188 17220 36430
rect 18956 27860 19012 27870
rect 18956 27766 19012 27804
rect 17164 27094 17220 27132
rect 17500 27746 17556 27758
rect 17500 27694 17502 27746
rect 17554 27694 17556 27746
rect 16716 26450 16772 26460
rect 17500 27076 17556 27694
rect 19516 27188 19572 37996
rect 19740 37986 19796 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 37156 20132 37166
rect 20188 37156 20244 41200
rect 20076 37154 20244 37156
rect 20076 37102 20078 37154
rect 20130 37102 20244 37154
rect 20076 37100 20244 37102
rect 20076 37090 20132 37100
rect 20860 36708 20916 41200
rect 21420 38052 21476 38062
rect 20860 36642 20916 36652
rect 20972 38050 21476 38052
rect 20972 37998 21422 38050
rect 21474 37998 21476 38050
rect 20972 37996 21476 37998
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 17612 27076 17668 27086
rect 17500 27074 17668 27076
rect 17500 27022 17614 27074
rect 17666 27022 17668 27074
rect 17500 27020 17668 27022
rect 16828 26292 16884 26302
rect 16828 26198 16884 26236
rect 16604 25508 16660 26124
rect 16604 25442 16660 25452
rect 17500 26178 17556 27020
rect 17612 27010 17668 27020
rect 18396 26962 18452 26974
rect 18396 26910 18398 26962
rect 18450 26910 18452 26962
rect 18396 26908 18452 26910
rect 18396 26852 18788 26908
rect 18508 26516 18564 26526
rect 17500 26126 17502 26178
rect 17554 26126 17556 26178
rect 16492 25330 16548 25340
rect 16268 25284 16324 25294
rect 16268 25190 16324 25228
rect 17500 25284 17556 26126
rect 17500 25218 17556 25228
rect 17612 26292 17668 26302
rect 17612 24946 17668 26236
rect 17612 24894 17614 24946
rect 17666 24894 17668 24946
rect 17612 24882 17668 24894
rect 18508 26290 18564 26460
rect 18732 26514 18788 26852
rect 18732 26462 18734 26514
rect 18786 26462 18788 26514
rect 18732 26450 18788 26462
rect 18844 26740 18900 26750
rect 18508 26238 18510 26290
rect 18562 26238 18564 26290
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 15932 24052 15988 24062
rect 15932 23958 15988 23996
rect 15148 23938 15540 23940
rect 15148 23886 15486 23938
rect 15538 23886 15540 23938
rect 15148 23884 15540 23886
rect 14812 23772 14980 23828
rect 14588 22484 14644 22494
rect 14588 22390 14644 22428
rect 14476 22306 14532 22316
rect 14140 22206 14142 22258
rect 14194 22206 14196 22258
rect 14140 22194 14196 22206
rect 14700 22148 14756 22158
rect 14700 22146 14868 22148
rect 14700 22094 14702 22146
rect 14754 22094 14868 22146
rect 14700 22092 14868 22094
rect 14700 22082 14756 22092
rect 12124 21746 12180 21756
rect 14700 21812 14756 21822
rect 14700 21718 14756 21756
rect 14812 21698 14868 22092
rect 14812 21646 14814 21698
rect 14866 21646 14868 21698
rect 14812 21634 14868 21646
rect 4172 21410 4228 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 14924 20188 14980 23772
rect 15036 22372 15092 22382
rect 15036 21586 15092 22316
rect 15036 21534 15038 21586
rect 15090 21534 15092 21586
rect 15036 21522 15092 21534
rect 14700 20132 14756 20142
rect 13916 20020 13972 20030
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1932 19346 1988 19358
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 18900 1988 19294
rect 4284 19236 4340 19246
rect 4284 19142 4340 19180
rect 11788 19124 11844 19134
rect 1932 18834 1988 18844
rect 9996 19012 10052 19022
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 9996 17778 10052 18956
rect 11116 18452 11172 18462
rect 11116 18358 11172 18396
rect 11788 18450 11844 19068
rect 11788 18398 11790 18450
rect 11842 18398 11844 18450
rect 11788 18386 11844 18398
rect 12796 18452 12852 18462
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 9996 17714 10052 17726
rect 12124 18228 12180 18238
rect 12124 17778 12180 18172
rect 12124 17726 12126 17778
rect 12178 17726 12180 17778
rect 12124 17714 12180 17726
rect 12796 17668 12852 18396
rect 13916 18338 13972 19964
rect 14700 19234 14756 20076
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14700 19170 14756 19182
rect 14812 20132 14980 20188
rect 15036 21140 15092 21150
rect 13916 18286 13918 18338
rect 13970 18286 13972 18338
rect 13916 18274 13972 18286
rect 14028 19010 14084 19022
rect 14028 18958 14030 19010
rect 14082 18958 14084 19010
rect 14028 18676 14084 18958
rect 14140 19010 14196 19022
rect 14140 18958 14142 19010
rect 14194 18958 14196 19010
rect 14140 18676 14196 18958
rect 14252 19012 14308 19022
rect 14252 18918 14308 18956
rect 14140 18620 14644 18676
rect 14028 18340 14084 18620
rect 14588 18562 14644 18620
rect 14588 18510 14590 18562
rect 14642 18510 14644 18562
rect 14588 18498 14644 18510
rect 14812 18450 14868 20132
rect 15036 19458 15092 21084
rect 15148 19684 15204 23884
rect 15484 23874 15540 23884
rect 16156 23938 16212 23950
rect 16156 23886 16158 23938
rect 16210 23886 16212 23938
rect 15708 23828 15764 23838
rect 15708 23734 15764 23772
rect 15596 23716 15652 23726
rect 15596 23622 15652 23660
rect 16156 23716 16212 23886
rect 16716 23940 16772 23950
rect 16492 23716 16548 23726
rect 16156 23714 16548 23716
rect 16156 23662 16494 23714
rect 16546 23662 16548 23714
rect 16156 23660 16548 23662
rect 15708 23156 15764 23166
rect 15596 22484 15652 22494
rect 15596 22370 15652 22428
rect 15596 22318 15598 22370
rect 15650 22318 15652 22370
rect 15484 21588 15540 21598
rect 15484 21494 15540 21532
rect 15260 21362 15316 21374
rect 15260 21310 15262 21362
rect 15314 21310 15316 21362
rect 15260 19908 15316 21310
rect 15484 20132 15540 20142
rect 15596 20132 15652 22318
rect 15708 22258 15764 23100
rect 15708 22206 15710 22258
rect 15762 22206 15764 22258
rect 15708 22194 15764 22206
rect 15820 23042 15876 23054
rect 15820 22990 15822 23042
rect 15874 22990 15876 23042
rect 15820 22148 15876 22990
rect 16156 22260 16212 23660
rect 16492 23650 16548 23660
rect 16492 23154 16548 23166
rect 16492 23102 16494 23154
rect 16546 23102 16548 23154
rect 16492 23044 16548 23102
rect 16492 22978 16548 22988
rect 16604 22372 16660 22410
rect 16604 22306 16660 22316
rect 16156 22166 16212 22204
rect 16380 22258 16436 22270
rect 16380 22206 16382 22258
rect 16434 22206 16436 22258
rect 15820 22082 15876 22092
rect 15932 22146 15988 22158
rect 15932 22094 15934 22146
rect 15986 22094 15988 22146
rect 15932 22036 15988 22094
rect 16380 22036 16436 22206
rect 16492 22148 16548 22158
rect 16492 22054 16548 22092
rect 15932 21980 16436 22036
rect 15820 21812 15876 21822
rect 15820 21586 15876 21756
rect 15820 21534 15822 21586
rect 15874 21534 15876 21586
rect 15820 21140 15876 21534
rect 15820 21074 15876 21084
rect 15540 20076 15652 20132
rect 16492 20132 16548 20142
rect 16716 20132 16772 23884
rect 17836 23940 17892 24670
rect 17836 23874 17892 23884
rect 17276 23828 17332 23838
rect 17276 23734 17332 23772
rect 17612 23492 17668 23502
rect 16940 23044 16996 23054
rect 16828 22370 16884 22382
rect 16828 22318 16830 22370
rect 16882 22318 16884 22370
rect 16828 21700 16884 22318
rect 16828 21634 16884 21644
rect 16940 20692 16996 22988
rect 17500 23044 17556 23054
rect 17500 22950 17556 22988
rect 17388 22482 17444 22494
rect 17388 22430 17390 22482
rect 17442 22430 17444 22482
rect 17388 22372 17444 22430
rect 17388 22306 17444 22316
rect 17612 22484 17668 23436
rect 17724 22596 17780 22606
rect 17724 22502 17780 22540
rect 18508 22596 18564 26238
rect 18844 26292 18900 26684
rect 19516 26628 19572 27132
rect 19628 27746 19684 27758
rect 19628 27694 19630 27746
rect 19682 27694 19684 27746
rect 19628 26852 19684 27694
rect 20524 27188 20580 27198
rect 20524 27094 20580 27132
rect 19628 26786 19684 26796
rect 20748 26852 20804 26862
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19516 26572 19684 26628
rect 19836 26618 20100 26628
rect 19628 26516 19684 26572
rect 19740 26516 19796 26526
rect 18844 26198 18900 26236
rect 19068 26460 19572 26516
rect 19628 26514 19796 26516
rect 19628 26462 19742 26514
rect 19794 26462 19796 26514
rect 19628 26460 19796 26462
rect 19068 25284 19124 26460
rect 19516 26402 19572 26460
rect 19740 26450 19796 26460
rect 20748 26514 20804 26796
rect 20748 26462 20750 26514
rect 20802 26462 20804 26514
rect 20748 26450 20804 26462
rect 19516 26350 19518 26402
rect 19570 26350 19572 26402
rect 19516 26338 19572 26350
rect 19964 26404 20020 26414
rect 19964 26310 20020 26348
rect 19180 26290 19236 26302
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 19180 26180 19236 26238
rect 19852 26292 19908 26302
rect 19628 26180 19684 26190
rect 19180 26178 19684 26180
rect 19180 26126 19630 26178
rect 19682 26126 19684 26178
rect 19180 26124 19684 26126
rect 19628 26114 19684 26124
rect 19852 25394 19908 26236
rect 20412 26292 20468 26302
rect 20412 26198 20468 26236
rect 20748 26292 20804 26302
rect 20748 26290 20916 26292
rect 20748 26238 20750 26290
rect 20802 26238 20916 26290
rect 20748 26236 20916 26238
rect 20748 26226 20804 26236
rect 19852 25342 19854 25394
rect 19906 25342 19908 25394
rect 19852 25330 19908 25342
rect 19068 23828 19124 25228
rect 20188 25282 20244 25294
rect 20188 25230 20190 25282
rect 20242 25230 20244 25282
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 25060 20244 25230
rect 20636 25284 20692 25294
rect 20636 25190 20692 25228
rect 20188 25004 20804 25060
rect 20748 24946 20804 25004
rect 20748 24894 20750 24946
rect 20802 24894 20804 24946
rect 19516 24050 19572 24062
rect 19516 23998 19518 24050
rect 19570 23998 19572 24050
rect 19068 23762 19124 23772
rect 19404 23828 19460 23838
rect 19404 23734 19460 23772
rect 19516 23268 19572 23998
rect 20636 23828 20692 23838
rect 19628 23714 19684 23726
rect 19628 23662 19630 23714
rect 19682 23662 19684 23714
rect 19628 23492 19684 23662
rect 19852 23716 19908 23754
rect 19852 23650 19908 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23426 19684 23436
rect 19516 23212 19908 23268
rect 18956 23156 19012 23166
rect 18956 23062 19012 23100
rect 18508 22530 18564 22540
rect 19628 23042 19684 23054
rect 19628 22990 19630 23042
rect 19682 22990 19684 23042
rect 17052 22260 17108 22270
rect 17500 22260 17556 22270
rect 17612 22260 17668 22428
rect 19628 22482 19684 22990
rect 19628 22430 19630 22482
rect 19682 22430 19684 22482
rect 19628 22418 19684 22430
rect 17052 22258 17220 22260
rect 17052 22206 17054 22258
rect 17106 22206 17220 22258
rect 17052 22204 17220 22206
rect 17052 22194 17108 22204
rect 17052 20692 17108 20702
rect 16940 20690 17108 20692
rect 16940 20638 17054 20690
rect 17106 20638 17108 20690
rect 16940 20636 17108 20638
rect 16492 20130 16772 20132
rect 16492 20078 16494 20130
rect 16546 20078 16772 20130
rect 16492 20076 16772 20078
rect 15484 20038 15540 20076
rect 15820 20020 15876 20030
rect 16156 20020 16212 20030
rect 15820 20018 15988 20020
rect 15820 19966 15822 20018
rect 15874 19966 15988 20018
rect 15820 19964 15988 19966
rect 15820 19954 15876 19964
rect 15260 19852 15764 19908
rect 15148 19628 15428 19684
rect 15036 19406 15038 19458
rect 15090 19406 15092 19458
rect 15036 19394 15092 19406
rect 15372 19460 15428 19628
rect 15708 19460 15764 19852
rect 15820 19460 15876 19470
rect 15372 19458 15540 19460
rect 15372 19406 15374 19458
rect 15426 19406 15540 19458
rect 15372 19404 15540 19406
rect 15708 19458 15876 19460
rect 15708 19406 15822 19458
rect 15874 19406 15876 19458
rect 15708 19404 15876 19406
rect 15372 19394 15428 19404
rect 15260 19348 15316 19358
rect 15148 19292 15260 19348
rect 14924 19124 14980 19134
rect 14924 19030 14980 19068
rect 14812 18398 14814 18450
rect 14866 18398 14868 18450
rect 14028 18284 14420 18340
rect 13916 17890 13972 17902
rect 13916 17838 13918 17890
rect 13970 17838 13972 17890
rect 12796 17574 12852 17612
rect 13580 17668 13636 17678
rect 4284 16882 4340 16894
rect 4284 16830 4286 16882
rect 4338 16830 4340 16882
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 1932 16146 1988 16156
rect 2044 16210 2100 16222
rect 2044 16158 2046 16210
rect 2098 16158 2100 16210
rect 2044 15540 2100 16158
rect 2044 15474 2100 15484
rect 4060 16098 4116 16110
rect 4060 16046 4062 16098
rect 4114 16046 4116 16098
rect 1932 15092 1988 15102
rect 1932 14998 1988 15036
rect 4060 14308 4116 16046
rect 4284 15764 4340 16830
rect 12796 16884 12852 16894
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4284 15698 4340 15708
rect 10668 15764 10724 15774
rect 4284 15428 4340 15438
rect 4284 15314 4340 15372
rect 4284 15262 4286 15314
rect 4338 15262 4340 15314
rect 4284 15250 4340 15262
rect 10668 15202 10724 15708
rect 12796 15426 12852 16828
rect 12796 15374 12798 15426
rect 12850 15374 12852 15426
rect 12796 15362 12852 15374
rect 13468 15874 13524 15886
rect 13468 15822 13470 15874
rect 13522 15822 13524 15874
rect 13468 15428 13524 15822
rect 13468 15362 13524 15372
rect 13580 15316 13636 17612
rect 13916 16994 13972 17838
rect 14140 17668 14196 17678
rect 14140 17574 14196 17612
rect 13916 16942 13918 16994
rect 13970 16942 13972 16994
rect 13916 16930 13972 16942
rect 14028 16884 14084 16894
rect 14028 16790 14084 16828
rect 14252 16882 14308 16894
rect 14252 16830 14254 16882
rect 14306 16830 14308 16882
rect 14252 16322 14308 16830
rect 14364 16770 14420 18284
rect 14700 18228 14756 18238
rect 14700 18134 14756 18172
rect 14588 17892 14644 17902
rect 14812 17892 14868 18398
rect 15148 18450 15204 19292
rect 15260 19254 15316 19292
rect 15148 18398 15150 18450
rect 15202 18398 15204 18450
rect 15148 18386 15204 18398
rect 15372 19012 15428 19022
rect 15372 18450 15428 18956
rect 15372 18398 15374 18450
rect 15426 18398 15428 18450
rect 15372 18386 15428 18398
rect 15484 18340 15540 19404
rect 15820 19394 15876 19404
rect 15932 19124 15988 19964
rect 16156 19926 16212 19964
rect 15932 19122 16100 19124
rect 15932 19070 15934 19122
rect 15986 19070 16100 19122
rect 15932 19068 16100 19070
rect 15932 19058 15988 19068
rect 15932 18452 15988 18462
rect 15932 18358 15988 18396
rect 15484 18274 15540 18284
rect 14588 17890 14868 17892
rect 14588 17838 14590 17890
rect 14642 17838 14868 17890
rect 14588 17836 14868 17838
rect 14588 17826 14644 17836
rect 14812 17554 14868 17836
rect 16044 17780 16100 19068
rect 16156 19122 16212 19134
rect 16156 19070 16158 19122
rect 16210 19070 16212 19122
rect 16156 18452 16212 19070
rect 16268 18564 16324 18574
rect 16268 18562 16436 18564
rect 16268 18510 16270 18562
rect 16322 18510 16436 18562
rect 16268 18508 16436 18510
rect 16268 18498 16324 18508
rect 16156 18340 16212 18396
rect 16380 18340 16436 18508
rect 16156 18284 16324 18340
rect 15484 17724 16100 17780
rect 15148 17668 15204 17678
rect 15484 17668 15540 17724
rect 15148 17666 15540 17668
rect 15148 17614 15150 17666
rect 15202 17614 15540 17666
rect 15148 17612 15540 17614
rect 16044 17668 16100 17724
rect 16268 17780 16324 18284
rect 16380 18116 16436 18284
rect 16492 18228 16548 20076
rect 16604 19348 16660 19358
rect 16604 19254 16660 19292
rect 16716 19236 16772 19246
rect 16716 19122 16772 19180
rect 16716 19070 16718 19122
rect 16770 19070 16772 19122
rect 16716 19058 16772 19070
rect 16940 19124 16996 19134
rect 16940 19030 16996 19068
rect 16492 18162 16548 18172
rect 16380 18050 16436 18060
rect 16268 17714 16324 17724
rect 16716 18004 16772 18014
rect 16156 17668 16212 17678
rect 16044 17666 16212 17668
rect 16044 17614 16158 17666
rect 16210 17614 16212 17666
rect 16044 17612 16212 17614
rect 15148 17602 15204 17612
rect 14812 17502 14814 17554
rect 14866 17502 14868 17554
rect 14812 17490 14868 17502
rect 15484 17554 15540 17612
rect 16156 17602 16212 17612
rect 16492 17668 16548 17678
rect 16492 17574 16548 17612
rect 16716 17666 16772 17948
rect 16716 17614 16718 17666
rect 16770 17614 16772 17666
rect 16716 17602 16772 17614
rect 15484 17502 15486 17554
rect 15538 17502 15540 17554
rect 15484 17490 15540 17502
rect 15820 17556 15876 17566
rect 15820 17462 15876 17500
rect 14700 17444 14756 17454
rect 14700 16882 14756 17388
rect 14700 16830 14702 16882
rect 14754 16830 14756 16882
rect 14700 16818 14756 16830
rect 15372 17444 15428 17454
rect 14364 16718 14366 16770
rect 14418 16718 14420 16770
rect 14364 16706 14420 16718
rect 14252 16270 14254 16322
rect 14306 16270 14308 16322
rect 14252 16258 14308 16270
rect 15260 16212 15316 16222
rect 14700 16210 15316 16212
rect 14700 16158 15262 16210
rect 15314 16158 15316 16210
rect 14700 16156 15316 16158
rect 13580 15222 13636 15260
rect 13692 16098 13748 16110
rect 13692 16046 13694 16098
rect 13746 16046 13748 16098
rect 13692 15988 13748 16046
rect 14140 15988 14196 15998
rect 13692 15986 14196 15988
rect 13692 15934 14142 15986
rect 14194 15934 14196 15986
rect 13692 15932 14196 15934
rect 13692 15764 13748 15932
rect 14140 15922 14196 15932
rect 10668 15150 10670 15202
rect 10722 15150 10724 15202
rect 10668 15138 10724 15150
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13692 14530 13748 15708
rect 14700 15426 14756 16156
rect 15260 16146 15316 16156
rect 15372 15986 15428 17388
rect 16492 17444 16548 17454
rect 16492 17350 16548 17388
rect 15596 16772 15652 16782
rect 15596 16322 15652 16716
rect 15596 16270 15598 16322
rect 15650 16270 15652 16322
rect 15596 16258 15652 16270
rect 15372 15934 15374 15986
rect 15426 15934 15428 15986
rect 15372 15922 15428 15934
rect 14700 15374 14702 15426
rect 14754 15374 14756 15426
rect 14700 15362 14756 15374
rect 13916 15316 13972 15326
rect 16940 15316 16996 15326
rect 17052 15316 17108 20636
rect 17164 17892 17220 22204
rect 17500 22258 17668 22260
rect 17500 22206 17502 22258
rect 17554 22206 17668 22258
rect 17500 22204 17668 22206
rect 19292 22370 19348 22382
rect 19292 22318 19294 22370
rect 19346 22318 19348 22370
rect 17500 22194 17556 22204
rect 18396 21812 18452 21822
rect 18396 21698 18452 21756
rect 19292 21812 19348 22318
rect 19852 22370 19908 23212
rect 19852 22318 19854 22370
rect 19906 22318 19908 22370
rect 19852 22306 19908 22318
rect 19516 22260 19572 22270
rect 19516 22166 19572 22204
rect 19740 22148 19796 22158
rect 19292 21746 19348 21756
rect 19628 22146 19796 22148
rect 19628 22094 19742 22146
rect 19794 22094 19796 22146
rect 19628 22092 19796 22094
rect 19628 21810 19684 22092
rect 19740 22082 19796 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21758 19630 21810
rect 19682 21758 19684 21810
rect 19628 21746 19684 21758
rect 19068 21700 19124 21710
rect 18396 21646 18398 21698
rect 18450 21646 18452 21698
rect 18060 21476 18116 21486
rect 18060 21382 18116 21420
rect 17836 20132 17892 20142
rect 17724 20076 17836 20132
rect 17612 20018 17668 20030
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 17612 19458 17668 19966
rect 17612 19406 17614 19458
rect 17666 19406 17668 19458
rect 17164 17668 17220 17836
rect 17164 17602 17220 17612
rect 17276 19124 17332 19134
rect 17276 18564 17332 19068
rect 17612 19124 17668 19406
rect 17612 19058 17668 19068
rect 17276 16772 17332 18508
rect 17388 19010 17444 19022
rect 17388 18958 17390 19010
rect 17442 18958 17444 19010
rect 17388 17668 17444 18958
rect 17500 19012 17556 19022
rect 17500 18918 17556 18956
rect 17724 18674 17780 20076
rect 17836 20038 17892 20076
rect 17948 20018 18004 20030
rect 18284 20020 18340 20030
rect 17948 19966 17950 20018
rect 18002 19966 18004 20018
rect 17948 19908 18004 19966
rect 17948 19842 18004 19852
rect 18060 19964 18284 20020
rect 17724 18622 17726 18674
rect 17778 18622 17780 18674
rect 17724 18610 17780 18622
rect 17948 19010 18004 19022
rect 17948 18958 17950 19010
rect 18002 18958 18004 19010
rect 17948 18676 18004 18958
rect 17948 18610 18004 18620
rect 18060 18562 18116 19964
rect 18284 19926 18340 19964
rect 18396 19908 18452 21646
rect 18844 21698 19124 21700
rect 18844 21646 19070 21698
rect 19122 21646 19124 21698
rect 18844 21644 19124 21646
rect 18620 21588 18676 21598
rect 18844 21588 18900 21644
rect 19068 21634 19124 21644
rect 19404 21700 19460 21710
rect 18620 21586 18900 21588
rect 18620 21534 18622 21586
rect 18674 21534 18900 21586
rect 18620 21532 18900 21534
rect 18508 20132 18564 20142
rect 18508 20038 18564 20076
rect 18396 19852 18564 19908
rect 18172 19796 18228 19806
rect 18172 19236 18228 19740
rect 18172 19142 18228 19180
rect 18508 19012 18564 19852
rect 18620 19906 18676 21532
rect 18956 21476 19012 21486
rect 19404 21476 19460 21644
rect 18956 20018 19012 21420
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 18956 19954 19012 19966
rect 19180 21420 19460 21476
rect 19852 21698 19908 21710
rect 19852 21646 19854 21698
rect 19906 21646 19908 21698
rect 19852 21588 19908 21646
rect 19964 21700 20020 21710
rect 19964 21606 20020 21644
rect 18620 19854 18622 19906
rect 18674 19854 18676 19906
rect 18620 19842 18676 19854
rect 18844 19908 18900 19918
rect 18732 19236 18788 19246
rect 18732 19142 18788 19180
rect 18844 19124 18900 19852
rect 19068 19236 19124 19246
rect 18956 19124 19012 19134
rect 18844 19122 19012 19124
rect 18844 19070 18958 19122
rect 19010 19070 19012 19122
rect 18844 19068 19012 19070
rect 18956 19058 19012 19068
rect 18508 18956 18900 19012
rect 18060 18510 18062 18562
rect 18114 18510 18116 18562
rect 18060 18498 18116 18510
rect 17612 18450 17668 18462
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18340 17668 18398
rect 18172 18452 18228 18462
rect 18172 18358 18228 18396
rect 18732 18450 18788 18462
rect 18732 18398 18734 18450
rect 18786 18398 18788 18450
rect 17388 17602 17444 17612
rect 17500 18284 17612 18340
rect 17500 17556 17556 18284
rect 17612 18274 17668 18284
rect 18732 18340 18788 18398
rect 18284 18228 18340 18238
rect 18508 18228 18564 18238
rect 17612 18116 17668 18126
rect 17612 17666 17668 18060
rect 17948 18116 18004 18126
rect 17948 17890 18004 18060
rect 17948 17838 17950 17890
rect 18002 17838 18004 17890
rect 17948 17826 18004 17838
rect 17612 17614 17614 17666
rect 17666 17614 17668 17666
rect 17612 17602 17668 17614
rect 18060 17668 18116 17678
rect 18060 17574 18116 17612
rect 17500 17490 17556 17500
rect 18284 17556 18340 18172
rect 18396 18172 18508 18228
rect 18396 17892 18452 18172
rect 18508 18162 18564 18172
rect 18396 17826 18452 17836
rect 17948 17442 18004 17454
rect 17948 17390 17950 17442
rect 18002 17390 18004 17442
rect 17612 17108 17668 17118
rect 17612 17014 17668 17052
rect 17388 16772 17444 16782
rect 17276 16770 17444 16772
rect 17276 16718 17390 16770
rect 17442 16718 17444 16770
rect 17276 16716 17444 16718
rect 17388 16706 17444 16716
rect 17500 16772 17556 16782
rect 17500 16678 17556 16716
rect 13972 15260 14308 15316
rect 13916 15222 13972 15260
rect 14252 14642 14308 15260
rect 16996 15260 17108 15316
rect 17500 15316 17556 15326
rect 16828 15204 16884 15242
rect 16828 15138 16884 15148
rect 14252 14590 14254 14642
rect 14306 14590 14308 14642
rect 14252 14578 14308 14590
rect 13692 14478 13694 14530
rect 13746 14478 13748 14530
rect 13692 14466 13748 14478
rect 4060 14242 4116 14252
rect 13468 14308 13524 14318
rect 13468 14214 13524 14252
rect 16828 13972 16884 13982
rect 16940 13972 16996 15260
rect 17500 15222 17556 15260
rect 17948 15148 18004 17390
rect 18284 16098 18340 17500
rect 18396 17554 18452 17566
rect 18396 17502 18398 17554
rect 18450 17502 18452 17554
rect 18396 17108 18452 17502
rect 18396 17042 18452 17052
rect 18620 17444 18676 17454
rect 18284 16046 18286 16098
rect 18338 16046 18340 16098
rect 18284 16034 18340 16046
rect 18620 16098 18676 17388
rect 18620 16046 18622 16098
rect 18674 16046 18676 16098
rect 18620 16034 18676 16046
rect 18732 16098 18788 18284
rect 18732 16046 18734 16098
rect 18786 16046 18788 16098
rect 17836 15092 18004 15148
rect 18396 15874 18452 15886
rect 18396 15822 18398 15874
rect 18450 15822 18452 15874
rect 18396 15428 18452 15822
rect 17836 14418 17892 15092
rect 18284 14532 18340 14542
rect 18396 14532 18452 15372
rect 18732 15204 18788 16046
rect 18844 16100 18900 18956
rect 19068 18452 19124 19180
rect 19068 18358 19124 18396
rect 19180 18116 19236 21420
rect 19852 20580 19908 21532
rect 20076 20804 20132 20814
rect 20636 20804 20692 23772
rect 20748 21924 20804 24894
rect 20860 23828 20916 26236
rect 20860 23762 20916 23772
rect 20972 22372 21028 37996
rect 21420 37986 21476 37996
rect 21532 37492 21588 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 23548 38276 23604 41200
rect 23548 38210 23604 38220
rect 21532 37426 21588 37436
rect 22764 37492 22820 37502
rect 22764 37398 22820 37436
rect 24220 37492 24276 41200
rect 24220 37426 24276 37436
rect 21196 37266 21252 37278
rect 21196 37214 21198 37266
rect 21250 37214 21252 37266
rect 21084 26964 21140 26974
rect 21084 26290 21140 26908
rect 21196 26628 21252 37214
rect 21868 37266 21924 37278
rect 21868 37214 21870 37266
rect 21922 37214 21924 37266
rect 21756 36482 21812 36494
rect 21756 36430 21758 36482
rect 21810 36430 21812 36482
rect 21756 27748 21812 36430
rect 21420 27746 21812 27748
rect 21420 27694 21758 27746
rect 21810 27694 21812 27746
rect 21420 27692 21812 27694
rect 21308 26962 21364 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 21308 26852 21364 26910
rect 21420 26962 21476 27692
rect 21756 27682 21812 27692
rect 21420 26910 21422 26962
rect 21474 26910 21476 26962
rect 21420 26898 21476 26910
rect 21644 26964 21700 26974
rect 21644 26870 21700 26908
rect 21308 26786 21364 26796
rect 21196 26572 21476 26628
rect 21308 26404 21364 26414
rect 21308 26310 21364 26348
rect 21084 26238 21086 26290
rect 21138 26238 21140 26290
rect 21084 26226 21140 26238
rect 21084 25284 21140 25294
rect 21084 24946 21140 25228
rect 21084 24894 21086 24946
rect 21138 24894 21140 24946
rect 21084 24882 21140 24894
rect 21420 23938 21476 26572
rect 21644 26404 21700 26414
rect 21644 26310 21700 26348
rect 21868 25172 21924 37214
rect 22316 36708 22372 36718
rect 22316 36614 22372 36652
rect 24892 36708 24948 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 24892 36642 24948 36652
rect 25004 38050 25060 38062
rect 25004 37998 25006 38050
rect 25058 37998 25060 38050
rect 22316 27860 22372 27870
rect 22204 27804 22316 27860
rect 22204 27076 22260 27804
rect 22316 27766 22372 27804
rect 25004 27186 25060 37998
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 25564 37266 25620 37278
rect 25564 37214 25566 37266
rect 25618 37214 25620 37266
rect 25004 27134 25006 27186
rect 25058 27134 25060 27186
rect 22204 26982 22260 27020
rect 23324 27076 23380 27086
rect 22876 26964 22932 26974
rect 22316 26962 22932 26964
rect 22316 26910 22878 26962
rect 22930 26910 22932 26962
rect 22316 26908 22932 26910
rect 22316 26514 22372 26908
rect 22876 26898 22932 26908
rect 22316 26462 22318 26514
rect 22370 26462 22372 26514
rect 22316 26450 22372 26462
rect 22428 26404 22484 26414
rect 22428 26310 22484 26348
rect 22204 26290 22260 26302
rect 22204 26238 22206 26290
rect 22258 26238 22260 26290
rect 21420 23886 21422 23938
rect 21474 23886 21476 23938
rect 21420 23716 21476 23886
rect 21644 25116 21924 25172
rect 21980 25284 22036 25294
rect 21644 23826 21700 25116
rect 21644 23774 21646 23826
rect 21698 23774 21700 23826
rect 21644 23762 21700 23774
rect 21420 23548 21476 23660
rect 21420 23492 21812 23548
rect 20972 22316 21364 22372
rect 21308 22148 21364 22316
rect 21420 22370 21476 23492
rect 21756 23042 21812 23492
rect 21756 22990 21758 23042
rect 21810 22990 21812 23042
rect 21756 22978 21812 22990
rect 21420 22318 21422 22370
rect 21474 22318 21476 22370
rect 21420 22306 21476 22318
rect 21644 22148 21700 22158
rect 21308 22146 21700 22148
rect 21308 22094 21646 22146
rect 21698 22094 21700 22146
rect 21308 22092 21700 22094
rect 21644 22082 21700 22092
rect 20748 21868 21252 21924
rect 21196 21588 21252 21868
rect 21532 21700 21588 21710
rect 21532 21698 21812 21700
rect 21532 21646 21534 21698
rect 21586 21646 21812 21698
rect 21532 21644 21812 21646
rect 21532 21634 21588 21644
rect 21196 21586 21364 21588
rect 21196 21534 21198 21586
rect 21250 21534 21364 21586
rect 21196 21532 21364 21534
rect 21196 21522 21252 21532
rect 21196 20804 21252 20814
rect 20636 20802 21252 20804
rect 20636 20750 21198 20802
rect 21250 20750 21252 20802
rect 20636 20748 21252 20750
rect 20076 20710 20132 20748
rect 21196 20738 21252 20748
rect 19852 20514 19908 20524
rect 20524 20580 20580 20590
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19292 20132 19348 20142
rect 19292 19348 19348 20076
rect 19292 19234 19348 19292
rect 20188 19348 20244 19358
rect 19292 19182 19294 19234
rect 19346 19182 19348 19234
rect 19292 19170 19348 19182
rect 19964 19236 20020 19246
rect 19964 19142 20020 19180
rect 20188 19234 20244 19292
rect 20188 19182 20190 19234
rect 20242 19182 20244 19234
rect 20188 19170 20244 19182
rect 19628 19124 19684 19134
rect 19628 19030 19684 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19292 18564 19348 18574
rect 19740 18564 19796 18574
rect 19292 18562 19796 18564
rect 19292 18510 19294 18562
rect 19346 18510 19742 18562
rect 19794 18510 19796 18562
rect 19292 18508 19796 18510
rect 19292 18498 19348 18508
rect 19292 18116 19348 18126
rect 19180 18060 19292 18116
rect 19292 18050 19348 18060
rect 19180 17666 19236 17678
rect 19180 17614 19182 17666
rect 19234 17614 19236 17666
rect 19180 17556 19236 17614
rect 19180 17490 19236 17500
rect 19404 16884 19460 18508
rect 19740 18498 19796 18508
rect 19964 18450 20020 18462
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19852 17780 19908 17790
rect 19852 17686 19908 17724
rect 19964 17668 20020 18398
rect 20524 18450 20580 20524
rect 21308 19684 21364 21532
rect 21532 20692 21588 20702
rect 21532 20690 21700 20692
rect 21532 20638 21534 20690
rect 21586 20638 21700 20690
rect 21532 20636 21700 20638
rect 21532 20626 21588 20636
rect 21420 20578 21476 20590
rect 21420 20526 21422 20578
rect 21474 20526 21476 20578
rect 21420 19908 21476 20526
rect 21420 19842 21476 19852
rect 21308 19628 21588 19684
rect 21420 19348 21476 19358
rect 20860 19346 21476 19348
rect 20860 19294 21422 19346
rect 21474 19294 21476 19346
rect 20860 19292 21476 19294
rect 20748 19236 20804 19246
rect 20748 19142 20804 19180
rect 20748 18564 20804 18574
rect 20860 18564 20916 19292
rect 21420 19282 21476 19292
rect 20748 18562 20916 18564
rect 20748 18510 20750 18562
rect 20802 18510 20916 18562
rect 20748 18508 20916 18510
rect 21308 19122 21364 19134
rect 21308 19070 21310 19122
rect 21362 19070 21364 19122
rect 20748 18498 20804 18508
rect 20524 18398 20526 18450
rect 20578 18398 20580 18450
rect 20524 18386 20580 18398
rect 20860 18340 20916 18350
rect 19964 17602 20020 17612
rect 20076 17892 20132 17902
rect 20076 17554 20132 17836
rect 20076 17502 20078 17554
rect 20130 17502 20132 17554
rect 20076 17490 20132 17502
rect 20300 17666 20356 17678
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 20300 17444 20356 17614
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20300 17220 20356 17388
rect 20300 17154 20356 17164
rect 20524 17668 20580 17678
rect 19740 17108 19796 17118
rect 20076 17108 20132 17118
rect 19796 17052 20020 17108
rect 19740 17042 19796 17052
rect 19404 16818 19460 16828
rect 19964 16994 20020 17052
rect 20076 17014 20132 17052
rect 20524 17106 20580 17612
rect 20524 17054 20526 17106
rect 20578 17054 20580 17106
rect 20524 17042 20580 17054
rect 20860 17106 20916 18284
rect 21308 17780 21364 19070
rect 21532 19124 21588 19628
rect 21532 19030 21588 19068
rect 21420 18450 21476 18462
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18116 21476 18398
rect 21420 18050 21476 18060
rect 21308 17714 21364 17724
rect 21420 17892 21476 17902
rect 20860 17054 20862 17106
rect 20914 17054 20916 17106
rect 19964 16942 19966 16994
rect 20018 16942 20020 16994
rect 19180 16100 19236 16110
rect 18844 16098 19236 16100
rect 18844 16046 19182 16098
rect 19234 16046 19236 16098
rect 18844 16044 19236 16046
rect 19180 16034 19236 16044
rect 19516 16100 19572 16110
rect 19740 16100 19796 16110
rect 19516 16098 19684 16100
rect 19516 16046 19518 16098
rect 19570 16046 19684 16098
rect 19516 16044 19684 16046
rect 19516 16034 19572 16044
rect 19180 15874 19236 15886
rect 19180 15822 19182 15874
rect 19234 15822 19236 15874
rect 19180 15148 19236 15822
rect 19628 15540 19684 16044
rect 19740 16006 19796 16044
rect 19964 16100 20020 16942
rect 20300 16996 20356 17006
rect 20300 16902 20356 16940
rect 20524 16884 20580 16894
rect 19964 16098 20356 16100
rect 19964 16046 19966 16098
rect 20018 16046 20356 16098
rect 19964 16044 20356 16046
rect 19964 16034 20020 16044
rect 20300 15986 20356 16044
rect 20300 15934 20302 15986
rect 20354 15934 20356 15986
rect 20300 15922 20356 15934
rect 20524 16098 20580 16828
rect 20524 16046 20526 16098
rect 20578 16046 20580 16098
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20412 15652 20468 15662
rect 19628 15484 20132 15540
rect 19516 15428 19572 15438
rect 19516 15334 19572 15372
rect 19628 15316 19684 15326
rect 19964 15316 20020 15326
rect 19628 15314 20020 15316
rect 19628 15262 19630 15314
rect 19682 15262 19966 15314
rect 20018 15262 20020 15314
rect 19628 15260 20020 15262
rect 19628 15250 19684 15260
rect 19964 15250 20020 15260
rect 18732 15138 18788 15148
rect 18284 14530 18452 14532
rect 18284 14478 18286 14530
rect 18338 14478 18452 14530
rect 18284 14476 18452 14478
rect 18844 15092 19236 15148
rect 20076 15202 20132 15484
rect 20412 15538 20468 15596
rect 20412 15486 20414 15538
rect 20466 15486 20468 15538
rect 20412 15474 20468 15486
rect 20076 15150 20078 15202
rect 20130 15150 20132 15202
rect 20076 15138 20132 15150
rect 20188 15314 20244 15326
rect 20188 15262 20190 15314
rect 20242 15262 20244 15314
rect 20188 15148 20244 15262
rect 20524 15314 20580 16046
rect 20860 16100 20916 17054
rect 21196 17668 21252 17678
rect 21196 17106 21252 17612
rect 21420 17554 21476 17836
rect 21420 17502 21422 17554
rect 21474 17502 21476 17554
rect 21420 17490 21476 17502
rect 21532 17780 21588 17790
rect 21644 17780 21700 20636
rect 21532 17778 21700 17780
rect 21532 17726 21534 17778
rect 21586 17726 21700 17778
rect 21532 17724 21700 17726
rect 21756 18004 21812 21644
rect 21980 20580 22036 25228
rect 22204 24052 22260 26238
rect 22876 26292 22932 26302
rect 22876 26198 22932 26236
rect 22092 22484 22148 22494
rect 22092 21698 22148 22428
rect 22204 21810 22260 23996
rect 23212 23940 23268 23950
rect 23324 23940 23380 27020
rect 24668 26852 24724 26862
rect 23660 26516 23716 26526
rect 23660 26422 23716 26460
rect 24332 26516 24388 26526
rect 24332 26422 24388 26460
rect 24668 26514 24724 26796
rect 25004 26628 25060 27134
rect 25228 36482 25284 36494
rect 25228 36430 25230 36482
rect 25282 36430 25284 36482
rect 25228 26852 25284 36430
rect 25228 26786 25284 26796
rect 25004 26572 25284 26628
rect 24668 26462 24670 26514
rect 24722 26462 24724 26514
rect 24668 26450 24724 26462
rect 25228 26516 25284 26572
rect 25228 26422 25284 26460
rect 25564 26514 25620 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 26124 36708 26180 36718
rect 26124 36614 26180 36652
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25676 27076 25732 27086
rect 25676 26982 25732 27020
rect 25564 26462 25566 26514
rect 25618 26462 25620 26514
rect 25564 26450 25620 26462
rect 23436 26292 23492 26302
rect 23772 26292 23828 26302
rect 23436 26198 23492 26236
rect 23660 26290 23828 26292
rect 23660 26238 23774 26290
rect 23826 26238 23828 26290
rect 23660 26236 23828 26238
rect 23212 23938 23380 23940
rect 23212 23886 23214 23938
rect 23266 23886 23380 23938
rect 23212 23884 23380 23886
rect 22428 23156 22484 23166
rect 22428 23062 22484 23100
rect 23212 23156 23268 23884
rect 23268 23100 23380 23156
rect 23212 23090 23268 23100
rect 22204 21758 22206 21810
rect 22258 21758 22260 21810
rect 22204 21746 22260 21758
rect 22316 22596 22372 22606
rect 22092 21646 22094 21698
rect 22146 21646 22148 21698
rect 22092 21634 22148 21646
rect 22204 20580 22260 20590
rect 21980 20578 22260 20580
rect 21980 20526 21982 20578
rect 22034 20526 22206 20578
rect 22258 20526 22260 20578
rect 21980 20524 22260 20526
rect 21980 20514 22036 20524
rect 22204 20514 22260 20524
rect 22316 19234 22372 22540
rect 22764 22484 22820 22494
rect 22652 20804 22708 20814
rect 22540 20578 22596 20590
rect 22540 20526 22542 20578
rect 22594 20526 22596 20578
rect 22540 19908 22596 20526
rect 22652 20130 22708 20748
rect 22652 20078 22654 20130
rect 22706 20078 22708 20130
rect 22652 20066 22708 20078
rect 22540 19852 22708 19908
rect 22316 19182 22318 19234
rect 22370 19182 22372 19234
rect 21980 18674 22036 18686
rect 21980 18622 21982 18674
rect 22034 18622 22036 18674
rect 21980 18452 22036 18622
rect 22316 18674 22372 19182
rect 22652 19122 22708 19852
rect 22652 19070 22654 19122
rect 22706 19070 22708 19122
rect 22540 19012 22596 19022
rect 22540 18918 22596 18956
rect 22316 18622 22318 18674
rect 22370 18622 22372 18674
rect 22316 18610 22372 18622
rect 21980 18386 22036 18396
rect 22316 18450 22372 18462
rect 22316 18398 22318 18450
rect 22370 18398 22372 18450
rect 21196 17054 21198 17106
rect 21250 17054 21252 17106
rect 21196 17042 21252 17054
rect 21420 17220 21476 17230
rect 21420 16882 21476 17164
rect 21532 17108 21588 17724
rect 21644 17556 21700 17566
rect 21756 17556 21812 17948
rect 22204 17556 22260 17566
rect 21644 17554 22204 17556
rect 21644 17502 21646 17554
rect 21698 17502 22204 17554
rect 21644 17500 22204 17502
rect 21644 17490 21700 17500
rect 21756 17220 21812 17230
rect 21812 17164 21924 17220
rect 21756 17154 21812 17164
rect 21532 17042 21588 17052
rect 21420 16830 21422 16882
rect 21474 16830 21476 16882
rect 21420 16818 21476 16830
rect 21868 16210 21924 17164
rect 22204 16996 22260 17500
rect 22316 17220 22372 18398
rect 22652 17780 22708 19070
rect 22764 18564 22820 22428
rect 23324 22372 23380 23100
rect 23324 22278 23380 22316
rect 23548 22930 23604 22942
rect 23548 22878 23550 22930
rect 23602 22878 23604 22930
rect 23324 22148 23380 22158
rect 22876 20580 22932 20590
rect 22876 19236 22932 20524
rect 23324 19236 23380 22092
rect 22876 19234 23044 19236
rect 22876 19182 22878 19234
rect 22930 19182 23044 19234
rect 22876 19180 23044 19182
rect 22876 19170 22932 19180
rect 22764 18562 22932 18564
rect 22764 18510 22766 18562
rect 22818 18510 22932 18562
rect 22764 18508 22932 18510
rect 22764 18498 22820 18508
rect 22652 17714 22708 17724
rect 22316 17154 22372 17164
rect 22316 16996 22372 17006
rect 22204 16994 22372 16996
rect 22204 16942 22318 16994
rect 22370 16942 22372 16994
rect 22204 16940 22372 16942
rect 22316 16930 22372 16940
rect 22540 16884 22596 16894
rect 21868 16158 21870 16210
rect 21922 16158 21924 16210
rect 21868 16146 21924 16158
rect 22428 16882 22596 16884
rect 22428 16830 22542 16882
rect 22594 16830 22596 16882
rect 22428 16828 22596 16830
rect 20860 16034 20916 16044
rect 22316 16100 22372 16110
rect 22428 16100 22484 16828
rect 22540 16818 22596 16828
rect 22316 16098 22484 16100
rect 22316 16046 22318 16098
rect 22370 16046 22484 16098
rect 22316 16044 22484 16046
rect 22316 15540 22372 16044
rect 22652 15876 22708 15886
rect 22316 15474 22372 15484
rect 22428 15874 22708 15876
rect 22428 15822 22654 15874
rect 22706 15822 22708 15874
rect 22428 15820 22708 15822
rect 22428 15652 22484 15820
rect 22652 15810 22708 15820
rect 22428 15538 22484 15596
rect 22428 15486 22430 15538
rect 22482 15486 22484 15538
rect 22428 15474 22484 15486
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 20524 15250 20580 15262
rect 22204 15314 22260 15326
rect 22204 15262 22206 15314
rect 22258 15262 22260 15314
rect 20188 15092 20916 15148
rect 18284 14466 18340 14476
rect 17836 14366 17838 14418
rect 17890 14366 17892 14418
rect 17836 14354 17892 14366
rect 18060 14306 18116 14318
rect 18060 14254 18062 14306
rect 18114 14254 18116 14306
rect 16828 13970 16996 13972
rect 16828 13918 16830 13970
rect 16882 13918 16996 13970
rect 16828 13916 16996 13918
rect 16828 13906 16884 13916
rect 16940 13412 16996 13916
rect 17612 13972 17668 13982
rect 18060 13972 18116 14254
rect 17612 13970 18116 13972
rect 17612 13918 17614 13970
rect 17666 13918 18116 13970
rect 17612 13916 18116 13918
rect 18172 14306 18228 14318
rect 18172 14254 18174 14306
rect 18226 14254 18228 14306
rect 17612 13906 17668 13916
rect 17948 13746 18004 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 16940 13346 16996 13356
rect 17500 13634 17556 13646
rect 17500 13582 17502 13634
rect 17554 13582 17556 13634
rect 4476 13290 4740 13300
rect 15820 13076 15876 13086
rect 15820 12982 15876 13020
rect 17500 13076 17556 13582
rect 17948 13412 18004 13694
rect 17948 13346 18004 13356
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17500 3556 17556 13020
rect 17948 13076 18004 13086
rect 18172 13076 18228 14254
rect 18732 13860 18788 13870
rect 18844 13860 18900 15092
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 18732 13858 18900 13860
rect 18732 13806 18734 13858
rect 18786 13806 18900 13858
rect 18732 13804 18900 13806
rect 18732 13794 18788 13804
rect 20860 13636 20916 15092
rect 21532 14532 21588 14542
rect 21980 14532 22036 14542
rect 21196 14530 22036 14532
rect 21196 14478 21534 14530
rect 21586 14478 21982 14530
rect 22034 14478 22036 14530
rect 21196 14476 22036 14478
rect 20860 13634 21028 13636
rect 20860 13582 20862 13634
rect 20914 13582 21028 13634
rect 20860 13580 21028 13582
rect 20860 13570 20916 13580
rect 17948 13074 18228 13076
rect 17948 13022 17950 13074
rect 18002 13022 18228 13074
rect 17948 13020 18228 13022
rect 18620 13412 18676 13422
rect 18620 13076 18676 13356
rect 19180 13076 19236 13086
rect 18620 13074 19236 13076
rect 18620 13022 19182 13074
rect 19234 13022 19236 13074
rect 18620 13020 19236 13022
rect 17948 13010 18004 13020
rect 18620 12962 18676 13020
rect 19180 13010 19236 13020
rect 18620 12910 18622 12962
rect 18674 12910 18676 12962
rect 18620 12898 18676 12910
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18620 3666 18676 3678
rect 18620 3614 18622 3666
rect 18674 3614 18676 3666
rect 17612 3556 17668 3566
rect 17500 3554 17668 3556
rect 17500 3502 17614 3554
rect 17666 3502 17668 3554
rect 17500 3500 17668 3502
rect 17612 3490 17668 3500
rect 18620 3388 18676 3614
rect 18172 3332 18676 3388
rect 20860 3668 20916 3678
rect 18172 800 18228 3332
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 3612
rect 20972 3556 21028 13580
rect 21196 13634 21252 14476
rect 21532 14466 21588 14476
rect 21980 14466 22036 14476
rect 21644 14308 21700 14318
rect 21644 14214 21700 14252
rect 22204 14308 22260 15262
rect 22876 15148 22932 18508
rect 22988 15986 23044 19180
rect 23324 19142 23380 19180
rect 23548 21364 23604 22878
rect 23660 22148 23716 26236
rect 23772 26226 23828 26236
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 26124 24050 26180 24062
rect 26124 23998 26126 24050
rect 26178 23998 26180 24050
rect 23996 23826 24052 23838
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 23996 23266 24052 23774
rect 23996 23214 23998 23266
rect 24050 23214 24052 23266
rect 23996 23202 24052 23214
rect 25340 23266 25396 23278
rect 25340 23214 25342 23266
rect 25394 23214 25396 23266
rect 24108 23154 24164 23166
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 23772 22932 23828 22942
rect 23772 22930 23940 22932
rect 23772 22878 23774 22930
rect 23826 22878 23940 22930
rect 23772 22876 23940 22878
rect 23772 22866 23828 22876
rect 23884 22260 23940 22876
rect 24108 22484 24164 23102
rect 25340 23156 25396 23214
rect 25900 23268 25956 23278
rect 26124 23268 26180 23998
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37884 23938 37940 23950
rect 37884 23886 37886 23938
rect 37938 23886 37940 23938
rect 25956 23212 26180 23268
rect 26572 23714 26628 23726
rect 26572 23662 26574 23714
rect 26626 23662 26628 23714
rect 25900 23174 25956 23212
rect 25340 23090 25396 23100
rect 25452 23156 25508 23166
rect 25788 23156 25844 23166
rect 25452 23154 25844 23156
rect 25452 23102 25454 23154
rect 25506 23102 25790 23154
rect 25842 23102 25844 23154
rect 25452 23100 25844 23102
rect 24332 23044 24388 23054
rect 24332 22950 24388 22988
rect 24108 22418 24164 22428
rect 24444 22932 24500 22942
rect 23772 22148 23828 22158
rect 23660 22092 23772 22148
rect 23772 22082 23828 22092
rect 23884 21586 23940 22204
rect 24108 22258 24164 22270
rect 24108 22206 24110 22258
rect 24162 22206 24164 22258
rect 24108 21698 24164 22206
rect 24108 21646 24110 21698
rect 24162 21646 24164 21698
rect 24108 21634 24164 21646
rect 24444 21698 24500 22876
rect 25340 22932 25396 22942
rect 25340 22838 25396 22876
rect 24444 21646 24446 21698
rect 24498 21646 24500 21698
rect 24444 21634 24500 21646
rect 25228 22372 25284 22382
rect 23884 21534 23886 21586
rect 23938 21534 23940 21586
rect 23884 21522 23940 21534
rect 24220 21586 24276 21598
rect 24220 21534 24222 21586
rect 24274 21534 24276 21586
rect 23660 21364 23716 21374
rect 23548 21362 23716 21364
rect 23548 21310 23662 21362
rect 23714 21310 23716 21362
rect 23548 21308 23716 21310
rect 23548 18900 23604 21308
rect 23660 21298 23716 21308
rect 24220 20188 24276 21534
rect 25228 20916 25284 22316
rect 25452 22148 25508 23100
rect 25788 23090 25844 23100
rect 26236 23156 26292 23166
rect 25900 23044 25956 23054
rect 25900 22930 25956 22988
rect 25900 22878 25902 22930
rect 25954 22878 25956 22930
rect 25900 22866 25956 22878
rect 26236 22484 26292 23100
rect 26236 22390 26292 22428
rect 26572 22372 26628 23662
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 37884 22484 37940 23886
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 37884 22418 37940 22428
rect 26684 22372 26740 22382
rect 26628 22370 26740 22372
rect 26628 22318 26686 22370
rect 26738 22318 26740 22370
rect 26628 22316 26740 22318
rect 26572 22306 26628 22316
rect 26684 22306 26740 22316
rect 25452 22082 25508 22092
rect 37884 21586 37940 21598
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 25228 20914 25732 20916
rect 25228 20862 25230 20914
rect 25282 20862 25732 20914
rect 25228 20860 25732 20862
rect 25228 20850 25284 20860
rect 23996 20132 24276 20188
rect 23548 18834 23604 18844
rect 23660 19010 23716 19022
rect 23660 18958 23662 19010
rect 23714 18958 23716 19010
rect 23212 18562 23268 18574
rect 23212 18510 23214 18562
rect 23266 18510 23268 18562
rect 23212 18228 23268 18510
rect 23548 18564 23604 18574
rect 23212 17668 23268 18172
rect 23436 18450 23492 18462
rect 23436 18398 23438 18450
rect 23490 18398 23492 18450
rect 23436 17892 23492 18398
rect 23212 17602 23268 17612
rect 23324 17836 23436 17892
rect 23324 16772 23380 17836
rect 23436 17826 23492 17836
rect 23548 17890 23604 18508
rect 23660 18340 23716 18958
rect 23660 18274 23716 18284
rect 23884 18228 23940 18238
rect 23996 18228 24052 20132
rect 24108 20020 24164 20030
rect 24108 19234 24164 19964
rect 24108 19182 24110 19234
rect 24162 19182 24164 19234
rect 24108 19170 24164 19182
rect 25676 20020 25732 20860
rect 29036 20020 29092 20030
rect 24780 19124 24836 19134
rect 24220 19122 24836 19124
rect 24220 19070 24782 19122
rect 24834 19070 24836 19122
rect 24220 19068 24836 19070
rect 24220 18674 24276 19068
rect 24780 19058 24836 19068
rect 24220 18622 24222 18674
rect 24274 18622 24276 18674
rect 24220 18610 24276 18622
rect 24332 18900 24388 18910
rect 24332 18674 24388 18844
rect 24332 18622 24334 18674
rect 24386 18622 24388 18674
rect 24332 18610 24388 18622
rect 24556 18676 24612 18686
rect 24556 18582 24612 18620
rect 24108 18564 24164 18574
rect 24108 18470 24164 18508
rect 24668 18564 24724 18574
rect 23940 18172 24052 18228
rect 24668 18228 24724 18508
rect 23884 18162 23940 18172
rect 23548 17838 23550 17890
rect 23602 17838 23604 17890
rect 23548 17826 23604 17838
rect 23548 17668 23604 17678
rect 23436 17556 23492 17566
rect 23436 17462 23492 17500
rect 23548 17554 23604 17612
rect 24668 17666 24724 18172
rect 25004 18564 25060 18574
rect 25004 17890 25060 18508
rect 25004 17838 25006 17890
rect 25058 17838 25060 17890
rect 25004 17826 25060 17838
rect 24668 17614 24670 17666
rect 24722 17614 24724 17666
rect 24668 17602 24724 17614
rect 25676 17666 25732 19964
rect 28588 19964 29036 20020
rect 26460 19908 26516 19918
rect 26124 19906 26516 19908
rect 26124 19854 26462 19906
rect 26514 19854 26516 19906
rect 26124 19852 26516 19854
rect 26012 19012 26068 19022
rect 26012 18674 26068 18956
rect 26012 18622 26014 18674
rect 26066 18622 26068 18674
rect 26012 18610 26068 18622
rect 26124 18674 26180 19852
rect 26460 19842 26516 19852
rect 27916 19908 27972 19918
rect 26908 19346 26964 19358
rect 26908 19294 26910 19346
rect 26962 19294 26964 19346
rect 26908 19236 26964 19294
rect 27916 19346 27972 19852
rect 28588 19906 28644 19964
rect 29036 19926 29092 19964
rect 37660 20018 37716 20030
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 29484 19908 29540 19918
rect 28588 19854 28590 19906
rect 28642 19854 28644 19906
rect 28588 19842 28644 19854
rect 29260 19852 29484 19908
rect 27916 19294 27918 19346
rect 27970 19294 27972 19346
rect 27916 19282 27972 19294
rect 28924 19794 28980 19806
rect 28924 19742 28926 19794
rect 28978 19742 28980 19794
rect 26908 19170 26964 19180
rect 27356 19236 27412 19246
rect 26124 18622 26126 18674
rect 26178 18622 26180 18674
rect 26124 18610 26180 18622
rect 26236 19124 26292 19134
rect 26236 18674 26292 19068
rect 27356 19122 27412 19180
rect 27356 19070 27358 19122
rect 27410 19070 27412 19122
rect 27356 19058 27412 19070
rect 27468 19122 27524 19134
rect 27468 19070 27470 19122
rect 27522 19070 27524 19122
rect 26236 18622 26238 18674
rect 26290 18622 26292 18674
rect 26236 18610 26292 18622
rect 27132 19010 27188 19022
rect 27132 18958 27134 19010
rect 27186 18958 27188 19010
rect 27132 18676 27188 18958
rect 27132 18610 27188 18620
rect 27020 18564 27076 18574
rect 27020 18470 27076 18508
rect 25788 18450 25844 18462
rect 25788 18398 25790 18450
rect 25842 18398 25844 18450
rect 25788 18228 25844 18398
rect 26348 18450 26404 18462
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 26124 18340 26180 18350
rect 26348 18340 26404 18398
rect 26796 18452 26852 18462
rect 26796 18358 26852 18396
rect 27244 18450 27300 18462
rect 27244 18398 27246 18450
rect 27298 18398 27300 18450
rect 26180 18284 26404 18340
rect 26460 18340 26516 18350
rect 26124 18274 26180 18284
rect 25788 18162 25844 18172
rect 26460 17778 26516 18284
rect 27132 18340 27188 18350
rect 27132 18246 27188 18284
rect 26460 17726 26462 17778
rect 26514 17726 26516 17778
rect 26460 17714 26516 17726
rect 27020 18228 27076 18238
rect 25676 17614 25678 17666
rect 25730 17614 25732 17666
rect 23548 17502 23550 17554
rect 23602 17502 23604 17554
rect 23548 17490 23604 17502
rect 24108 17556 24164 17566
rect 24108 17462 24164 17500
rect 24444 17554 24500 17566
rect 24444 17502 24446 17554
rect 24498 17502 24500 17554
rect 23324 16716 23604 16772
rect 22988 15934 22990 15986
rect 23042 15934 23044 15986
rect 22988 15922 23044 15934
rect 23324 15540 23380 15550
rect 23324 15314 23380 15484
rect 23324 15262 23326 15314
rect 23378 15262 23380 15314
rect 23324 15148 23380 15262
rect 23548 15316 23604 16716
rect 24220 16098 24276 16110
rect 24220 16046 24222 16098
rect 24274 16046 24276 16098
rect 24220 15426 24276 16046
rect 24220 15374 24222 15426
rect 24274 15374 24276 15426
rect 24220 15362 24276 15374
rect 24444 15986 24500 17502
rect 24892 17556 24948 17566
rect 24892 17462 24948 17500
rect 24444 15934 24446 15986
rect 24498 15934 24500 15986
rect 23548 15222 23604 15260
rect 22316 15092 22372 15102
rect 22316 14418 22372 15036
rect 22540 15092 22596 15102
rect 22876 15092 23156 15148
rect 23324 15092 23604 15148
rect 22540 14998 22596 15036
rect 23100 14644 23156 15092
rect 23100 14642 23380 14644
rect 23100 14590 23102 14642
rect 23154 14590 23380 14642
rect 23100 14588 23380 14590
rect 23100 14578 23156 14588
rect 22316 14366 22318 14418
rect 22370 14366 22372 14418
rect 22316 14354 22372 14366
rect 22204 14242 22260 14252
rect 22652 14308 22708 14318
rect 22652 14214 22708 14252
rect 23324 13858 23380 14588
rect 23548 14642 23604 15092
rect 24444 14756 24500 15934
rect 25676 16098 25732 17614
rect 27020 17332 27076 18172
rect 27244 17668 27300 18398
rect 27356 18452 27412 18462
rect 27468 18452 27524 19070
rect 28924 19124 28980 19742
rect 28924 19058 28980 19068
rect 27356 18450 27524 18452
rect 27356 18398 27358 18450
rect 27410 18398 27524 18450
rect 27356 18396 27524 18398
rect 27356 18228 27412 18396
rect 27356 18162 27412 18172
rect 28588 17778 28644 17790
rect 28588 17726 28590 17778
rect 28642 17726 28644 17778
rect 27804 17668 27860 17678
rect 27244 17612 27748 17668
rect 27020 17276 27412 17332
rect 26684 16996 26740 17006
rect 26684 16902 26740 16940
rect 27244 16994 27300 17006
rect 27244 16942 27246 16994
rect 27298 16942 27300 16994
rect 26460 16882 26516 16894
rect 26460 16830 26462 16882
rect 26514 16830 26516 16882
rect 26460 16210 26516 16830
rect 26796 16884 26852 16894
rect 27020 16884 27076 16894
rect 26796 16882 27076 16884
rect 26796 16830 26798 16882
rect 26850 16830 27022 16882
rect 27074 16830 27076 16882
rect 26796 16828 27076 16830
rect 26796 16818 26852 16828
rect 27020 16818 27076 16828
rect 27244 16884 27300 16942
rect 27356 16994 27412 17276
rect 27692 17106 27748 17612
rect 27692 17054 27694 17106
rect 27746 17054 27748 17106
rect 27692 17042 27748 17054
rect 27356 16942 27358 16994
rect 27410 16942 27412 16994
rect 27356 16930 27412 16942
rect 27804 16994 27860 17612
rect 28588 17668 28644 17726
rect 28588 17602 28644 17612
rect 29260 17778 29316 19852
rect 29484 19814 29540 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 19236 37716 19966
rect 37884 20020 37940 21534
rect 40012 21362 40068 21374
rect 40012 21310 40014 21362
rect 40066 21310 40068 21362
rect 40012 20916 40068 21310
rect 40012 20850 40068 20860
rect 37884 19954 37940 19964
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37660 19170 37716 19180
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 29260 17726 29262 17778
rect 29314 17726 29316 17778
rect 27804 16942 27806 16994
rect 27858 16942 27860 16994
rect 27804 16930 27860 16942
rect 27244 16818 27300 16828
rect 28588 16884 28644 16894
rect 26460 16158 26462 16210
rect 26514 16158 26516 16210
rect 26460 16146 26516 16158
rect 28588 16210 28644 16828
rect 28588 16158 28590 16210
rect 28642 16158 28644 16210
rect 28588 16146 28644 16158
rect 29260 16210 29316 17726
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 37660 16884 37716 16894
rect 37660 16790 37716 16828
rect 40012 16884 40068 16894
rect 40012 16770 40068 16828
rect 40012 16718 40014 16770
rect 40066 16718 40068 16770
rect 40012 16706 40068 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 29260 16158 29262 16210
rect 29314 16158 29316 16210
rect 29260 16146 29316 16158
rect 25676 16046 25678 16098
rect 25730 16046 25732 16098
rect 24444 14690 24500 14700
rect 25564 14756 25620 14766
rect 23548 14590 23550 14642
rect 23602 14590 23604 14642
rect 23548 14578 23604 14590
rect 24556 14644 24612 14654
rect 23324 13806 23326 13858
rect 23378 13806 23380 13858
rect 23324 13794 23380 13806
rect 24108 13748 24164 13758
rect 24556 13748 24612 14588
rect 25564 14420 25620 14700
rect 25676 14644 25732 16046
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 25676 14578 25732 14588
rect 26348 14644 26404 14654
rect 26348 14530 26404 14588
rect 26908 14644 26964 14654
rect 26908 14550 26964 14588
rect 26348 14478 26350 14530
rect 26402 14478 26404 14530
rect 26348 14466 26404 14478
rect 25676 14420 25732 14430
rect 25564 14418 25732 14420
rect 25564 14366 25678 14418
rect 25730 14366 25732 14418
rect 25564 14364 25732 14366
rect 25676 14354 25732 14364
rect 24108 13746 24612 13748
rect 24108 13694 24110 13746
rect 24162 13694 24558 13746
rect 24610 13694 24612 13746
rect 24108 13692 24612 13694
rect 24108 13682 24164 13692
rect 24556 13682 24612 13692
rect 21196 13582 21198 13634
rect 21250 13582 21252 13634
rect 21196 13570 21252 13582
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 21084 3556 21140 3566
rect 20972 3554 21140 3556
rect 20972 3502 21086 3554
rect 21138 3502 21140 3554
rect 20972 3500 21140 3502
rect 21084 3490 21140 3500
rect 18144 0 18256 800
rect 20832 0 20944 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 15372 38274 15428 38276
rect 15372 38222 15374 38274
rect 15374 38222 15426 38274
rect 15426 38222 15428 38274
rect 15372 38220 15428 38222
rect 16156 38220 16212 38276
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 16828 36652 16884 36708
rect 18060 36706 18116 36708
rect 18060 36654 18062 36706
rect 18062 36654 18114 36706
rect 18114 36654 18116 36706
rect 18060 36652 18116 36654
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 13804 28028 13860 28084
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 27074 4340 27076
rect 4284 27022 4286 27074
rect 4286 27022 4338 27074
rect 4338 27022 4340 27074
rect 4284 27020 4340 27022
rect 11228 27020 11284 27076
rect 1932 26236 1988 26292
rect 4172 26908 4228 26964
rect 1932 23548 1988 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 1932 22482 1988 22484
rect 1932 22430 1934 22482
rect 1934 22430 1986 22482
rect 1986 22430 1988 22482
rect 1932 22428 1988 22430
rect 13132 26796 13188 26852
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 14812 28082 14868 28084
rect 14812 28030 14814 28082
rect 14814 28030 14866 28082
rect 14866 28030 14868 28082
rect 14812 28028 14868 28030
rect 15036 27858 15092 27860
rect 15036 27806 15038 27858
rect 15038 27806 15090 27858
rect 15090 27806 15092 27858
rect 15036 27804 15092 27806
rect 14140 27020 14196 27076
rect 15036 27580 15092 27636
rect 14252 26908 14308 26964
rect 13356 25676 13412 25732
rect 14140 25394 14196 25396
rect 14140 25342 14142 25394
rect 14142 25342 14194 25394
rect 14194 25342 14196 25394
rect 14140 25340 14196 25342
rect 14812 25730 14868 25732
rect 14812 25678 14814 25730
rect 14814 25678 14866 25730
rect 14866 25678 14868 25730
rect 14812 25676 14868 25678
rect 15148 25676 15204 25732
rect 15596 26796 15652 26852
rect 16044 27858 16100 27860
rect 16044 27806 16046 27858
rect 16046 27806 16098 27858
rect 16098 27806 16100 27858
rect 16044 27804 16100 27806
rect 16044 27634 16100 27636
rect 16044 27582 16046 27634
rect 16046 27582 16098 27634
rect 16098 27582 16100 27634
rect 16044 27580 16100 27582
rect 16156 26684 16212 26740
rect 16268 27132 16324 27188
rect 16604 26796 16660 26852
rect 15372 25564 15428 25620
rect 15148 25452 15204 25508
rect 14812 25340 14868 25396
rect 13132 25228 13188 25284
rect 14364 25228 14420 25284
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 11004 23772 11060 23828
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 13692 23100 13748 23156
rect 13132 22540 13188 22596
rect 13580 22988 13636 23044
rect 9996 22482 10052 22484
rect 9996 22430 9998 22482
rect 9998 22430 10050 22482
rect 10050 22430 10052 22482
rect 9996 22428 10052 22430
rect 14364 23826 14420 23828
rect 14364 23774 14366 23826
rect 14366 23774 14418 23826
rect 14418 23774 14420 23826
rect 14364 23772 14420 23774
rect 13916 22988 13972 23044
rect 4284 22370 4340 22372
rect 4284 22318 4286 22370
rect 4286 22318 4338 22370
rect 4338 22318 4340 22370
rect 4284 22316 4340 22318
rect 12908 22370 12964 22372
rect 12908 22318 12910 22370
rect 12910 22318 12962 22370
rect 12962 22318 12964 22370
rect 12908 22316 12964 22318
rect 13580 22316 13636 22372
rect 13916 22540 13972 22596
rect 14252 23660 14308 23716
rect 14924 23996 14980 24052
rect 18956 27858 19012 27860
rect 18956 27806 18958 27858
rect 18958 27806 19010 27858
rect 19010 27806 19012 27858
rect 18956 27804 19012 27806
rect 17164 27186 17220 27188
rect 17164 27134 17166 27186
rect 17166 27134 17218 27186
rect 17218 27134 17220 27186
rect 17164 27132 17220 27134
rect 16716 26460 16772 26516
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20860 36652 20916 36708
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19516 27132 19572 27188
rect 16828 26290 16884 26292
rect 16828 26238 16830 26290
rect 16830 26238 16882 26290
rect 16882 26238 16884 26290
rect 16828 26236 16884 26238
rect 16604 26124 16660 26180
rect 16604 25452 16660 25508
rect 18508 26460 18564 26516
rect 16492 25340 16548 25396
rect 16268 25282 16324 25284
rect 16268 25230 16270 25282
rect 16270 25230 16322 25282
rect 16322 25230 16324 25282
rect 16268 25228 16324 25230
rect 17500 25228 17556 25284
rect 17612 26236 17668 26292
rect 18844 26684 18900 26740
rect 15932 24050 15988 24052
rect 15932 23998 15934 24050
rect 15934 23998 15986 24050
rect 15986 23998 15988 24050
rect 15932 23996 15988 23998
rect 14588 22482 14644 22484
rect 14588 22430 14590 22482
rect 14590 22430 14642 22482
rect 14642 22430 14644 22482
rect 14588 22428 14644 22430
rect 14476 22316 14532 22372
rect 12124 21756 12180 21812
rect 14700 21810 14756 21812
rect 14700 21758 14702 21810
rect 14702 21758 14754 21810
rect 14754 21758 14756 21810
rect 14700 21756 14756 21758
rect 4172 21420 4228 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 15036 22316 15092 22372
rect 14700 20076 14756 20132
rect 13916 19964 13972 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4284 19234 4340 19236
rect 4284 19182 4286 19234
rect 4286 19182 4338 19234
rect 4338 19182 4340 19234
rect 4284 19180 4340 19182
rect 11788 19068 11844 19124
rect 1932 18844 1988 18900
rect 9996 18956 10052 19012
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 11116 18450 11172 18452
rect 11116 18398 11118 18450
rect 11118 18398 11170 18450
rect 11170 18398 11172 18450
rect 11116 18396 11172 18398
rect 12796 18396 12852 18452
rect 12124 18172 12180 18228
rect 15036 21084 15092 21140
rect 14028 18620 14084 18676
rect 14252 19010 14308 19012
rect 14252 18958 14254 19010
rect 14254 18958 14306 19010
rect 14306 18958 14308 19010
rect 14252 18956 14308 18958
rect 15708 23826 15764 23828
rect 15708 23774 15710 23826
rect 15710 23774 15762 23826
rect 15762 23774 15764 23826
rect 15708 23772 15764 23774
rect 15596 23714 15652 23716
rect 15596 23662 15598 23714
rect 15598 23662 15650 23714
rect 15650 23662 15652 23714
rect 15596 23660 15652 23662
rect 16716 23938 16772 23940
rect 16716 23886 16718 23938
rect 16718 23886 16770 23938
rect 16770 23886 16772 23938
rect 16716 23884 16772 23886
rect 15708 23100 15764 23156
rect 15596 22428 15652 22484
rect 15484 21586 15540 21588
rect 15484 21534 15486 21586
rect 15486 21534 15538 21586
rect 15538 21534 15540 21586
rect 15484 21532 15540 21534
rect 16492 22988 16548 23044
rect 16604 22370 16660 22372
rect 16604 22318 16606 22370
rect 16606 22318 16658 22370
rect 16658 22318 16660 22370
rect 16604 22316 16660 22318
rect 16156 22258 16212 22260
rect 16156 22206 16158 22258
rect 16158 22206 16210 22258
rect 16210 22206 16212 22258
rect 16156 22204 16212 22206
rect 15820 22092 15876 22148
rect 16492 22146 16548 22148
rect 16492 22094 16494 22146
rect 16494 22094 16546 22146
rect 16546 22094 16548 22146
rect 16492 22092 16548 22094
rect 15820 21756 15876 21812
rect 15820 21084 15876 21140
rect 15484 20130 15540 20132
rect 15484 20078 15486 20130
rect 15486 20078 15538 20130
rect 15538 20078 15540 20130
rect 15484 20076 15540 20078
rect 17836 23884 17892 23940
rect 17276 23826 17332 23828
rect 17276 23774 17278 23826
rect 17278 23774 17330 23826
rect 17330 23774 17332 23826
rect 17276 23772 17332 23774
rect 17612 23436 17668 23492
rect 16940 22988 16996 23044
rect 16828 21644 16884 21700
rect 17500 23042 17556 23044
rect 17500 22990 17502 23042
rect 17502 22990 17554 23042
rect 17554 22990 17556 23042
rect 17500 22988 17556 22990
rect 17388 22316 17444 22372
rect 17724 22594 17780 22596
rect 17724 22542 17726 22594
rect 17726 22542 17778 22594
rect 17778 22542 17780 22594
rect 17724 22540 17780 22542
rect 20524 27186 20580 27188
rect 20524 27134 20526 27186
rect 20526 27134 20578 27186
rect 20578 27134 20580 27186
rect 20524 27132 20580 27134
rect 19628 26796 19684 26852
rect 20748 26796 20804 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 18844 26290 18900 26292
rect 18844 26238 18846 26290
rect 18846 26238 18898 26290
rect 18898 26238 18900 26290
rect 18844 26236 18900 26238
rect 19964 26402 20020 26404
rect 19964 26350 19966 26402
rect 19966 26350 20018 26402
rect 20018 26350 20020 26402
rect 19964 26348 20020 26350
rect 19852 26236 19908 26292
rect 20412 26290 20468 26292
rect 20412 26238 20414 26290
rect 20414 26238 20466 26290
rect 20466 26238 20468 26290
rect 20412 26236 20468 26238
rect 19068 25228 19124 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20636 25282 20692 25284
rect 20636 25230 20638 25282
rect 20638 25230 20690 25282
rect 20690 25230 20692 25282
rect 20636 25228 20692 25230
rect 19068 23772 19124 23828
rect 19404 23826 19460 23828
rect 19404 23774 19406 23826
rect 19406 23774 19458 23826
rect 19458 23774 19460 23826
rect 19404 23772 19460 23774
rect 20636 23772 20692 23828
rect 19852 23714 19908 23716
rect 19852 23662 19854 23714
rect 19854 23662 19906 23714
rect 19906 23662 19908 23714
rect 19852 23660 19908 23662
rect 19628 23436 19684 23492
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18956 23154 19012 23156
rect 18956 23102 18958 23154
rect 18958 23102 19010 23154
rect 19010 23102 19012 23154
rect 18956 23100 19012 23102
rect 18508 22540 18564 22596
rect 17612 22428 17668 22484
rect 15260 19346 15316 19348
rect 15260 19294 15262 19346
rect 15262 19294 15314 19346
rect 15314 19294 15316 19346
rect 15260 19292 15316 19294
rect 14924 19122 14980 19124
rect 14924 19070 14926 19122
rect 14926 19070 14978 19122
rect 14978 19070 14980 19122
rect 14924 19068 14980 19070
rect 12796 17666 12852 17668
rect 12796 17614 12798 17666
rect 12798 17614 12850 17666
rect 12850 17614 12852 17666
rect 12796 17612 12852 17614
rect 13580 17666 13636 17668
rect 13580 17614 13582 17666
rect 13582 17614 13634 17666
rect 13634 17614 13636 17666
rect 13580 17612 13636 17614
rect 1932 16156 1988 16212
rect 2044 15484 2100 15540
rect 1932 15090 1988 15092
rect 1932 15038 1934 15090
rect 1934 15038 1986 15090
rect 1986 15038 1988 15090
rect 1932 15036 1988 15038
rect 12796 16828 12852 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4284 15708 4340 15764
rect 10668 15708 10724 15764
rect 4284 15372 4340 15428
rect 13468 15372 13524 15428
rect 14140 17666 14196 17668
rect 14140 17614 14142 17666
rect 14142 17614 14194 17666
rect 14194 17614 14196 17666
rect 14140 17612 14196 17614
rect 14028 16882 14084 16884
rect 14028 16830 14030 16882
rect 14030 16830 14082 16882
rect 14082 16830 14084 16882
rect 14028 16828 14084 16830
rect 14700 18226 14756 18228
rect 14700 18174 14702 18226
rect 14702 18174 14754 18226
rect 14754 18174 14756 18226
rect 14700 18172 14756 18174
rect 15372 18956 15428 19012
rect 16156 20018 16212 20020
rect 16156 19966 16158 20018
rect 16158 19966 16210 20018
rect 16210 19966 16212 20018
rect 16156 19964 16212 19966
rect 15932 18450 15988 18452
rect 15932 18398 15934 18450
rect 15934 18398 15986 18450
rect 15986 18398 15988 18450
rect 15932 18396 15988 18398
rect 15484 18284 15540 18340
rect 16156 18396 16212 18452
rect 16380 18284 16436 18340
rect 16604 19346 16660 19348
rect 16604 19294 16606 19346
rect 16606 19294 16658 19346
rect 16658 19294 16660 19346
rect 16604 19292 16660 19294
rect 16716 19180 16772 19236
rect 16940 19122 16996 19124
rect 16940 19070 16942 19122
rect 16942 19070 16994 19122
rect 16994 19070 16996 19122
rect 16940 19068 16996 19070
rect 16492 18172 16548 18228
rect 16380 18060 16436 18116
rect 16268 17724 16324 17780
rect 16716 17948 16772 18004
rect 16492 17666 16548 17668
rect 16492 17614 16494 17666
rect 16494 17614 16546 17666
rect 16546 17614 16548 17666
rect 16492 17612 16548 17614
rect 15820 17554 15876 17556
rect 15820 17502 15822 17554
rect 15822 17502 15874 17554
rect 15874 17502 15876 17554
rect 15820 17500 15876 17502
rect 14700 17388 14756 17444
rect 15372 17388 15428 17444
rect 13580 15314 13636 15316
rect 13580 15262 13582 15314
rect 13582 15262 13634 15314
rect 13634 15262 13636 15314
rect 13580 15260 13636 15262
rect 13692 15708 13748 15764
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 16492 17442 16548 17444
rect 16492 17390 16494 17442
rect 16494 17390 16546 17442
rect 16546 17390 16548 17442
rect 16492 17388 16548 17390
rect 15596 16716 15652 16772
rect 18396 21756 18452 21812
rect 19516 22258 19572 22260
rect 19516 22206 19518 22258
rect 19518 22206 19570 22258
rect 19570 22206 19572 22258
rect 19516 22204 19572 22206
rect 19292 21756 19348 21812
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 18060 21474 18116 21476
rect 18060 21422 18062 21474
rect 18062 21422 18114 21474
rect 18114 21422 18116 21474
rect 18060 21420 18116 21422
rect 17836 20130 17892 20132
rect 17836 20078 17838 20130
rect 17838 20078 17890 20130
rect 17890 20078 17892 20130
rect 17836 20076 17892 20078
rect 17164 17836 17220 17892
rect 17164 17612 17220 17668
rect 17276 19068 17332 19124
rect 17612 19068 17668 19124
rect 17276 18508 17332 18564
rect 17500 19010 17556 19012
rect 17500 18958 17502 19010
rect 17502 18958 17554 19010
rect 17554 18958 17556 19010
rect 17500 18956 17556 18958
rect 17948 19852 18004 19908
rect 18284 20018 18340 20020
rect 18284 19966 18286 20018
rect 18286 19966 18338 20018
rect 18338 19966 18340 20018
rect 18284 19964 18340 19966
rect 17948 18620 18004 18676
rect 19404 21698 19460 21700
rect 19404 21646 19406 21698
rect 19406 21646 19458 21698
rect 19458 21646 19460 21698
rect 19404 21644 19460 21646
rect 18508 20130 18564 20132
rect 18508 20078 18510 20130
rect 18510 20078 18562 20130
rect 18562 20078 18564 20130
rect 18508 20076 18564 20078
rect 18172 19740 18228 19796
rect 18172 19234 18228 19236
rect 18172 19182 18174 19234
rect 18174 19182 18226 19234
rect 18226 19182 18228 19234
rect 18172 19180 18228 19182
rect 18956 21420 19012 21476
rect 19964 21698 20020 21700
rect 19964 21646 19966 21698
rect 19966 21646 20018 21698
rect 20018 21646 20020 21698
rect 19964 21644 20020 21646
rect 19852 21532 19908 21588
rect 18844 19852 18900 19908
rect 18732 19234 18788 19236
rect 18732 19182 18734 19234
rect 18734 19182 18786 19234
rect 18786 19182 18788 19234
rect 18732 19180 18788 19182
rect 19068 19180 19124 19236
rect 18172 18450 18228 18452
rect 18172 18398 18174 18450
rect 18174 18398 18226 18450
rect 18226 18398 18228 18450
rect 18172 18396 18228 18398
rect 17388 17612 17444 17668
rect 17612 18284 17668 18340
rect 18732 18284 18788 18340
rect 18284 18172 18340 18228
rect 17612 18060 17668 18116
rect 17948 18060 18004 18116
rect 18060 17666 18116 17668
rect 18060 17614 18062 17666
rect 18062 17614 18114 17666
rect 18114 17614 18116 17666
rect 18060 17612 18116 17614
rect 17500 17500 17556 17556
rect 18508 18172 18564 18228
rect 18396 17836 18452 17892
rect 18284 17500 18340 17556
rect 17612 17106 17668 17108
rect 17612 17054 17614 17106
rect 17614 17054 17666 17106
rect 17666 17054 17668 17106
rect 17612 17052 17668 17054
rect 17500 16770 17556 16772
rect 17500 16718 17502 16770
rect 17502 16718 17554 16770
rect 17554 16718 17556 16770
rect 17500 16716 17556 16718
rect 13916 15314 13972 15316
rect 13916 15262 13918 15314
rect 13918 15262 13970 15314
rect 13970 15262 13972 15314
rect 13916 15260 13972 15262
rect 16940 15260 16996 15316
rect 17500 15314 17556 15316
rect 17500 15262 17502 15314
rect 17502 15262 17554 15314
rect 17554 15262 17556 15314
rect 17500 15260 17556 15262
rect 16828 15202 16884 15204
rect 16828 15150 16830 15202
rect 16830 15150 16882 15202
rect 16882 15150 16884 15202
rect 16828 15148 16884 15150
rect 4060 14252 4116 14308
rect 13468 14306 13524 14308
rect 13468 14254 13470 14306
rect 13470 14254 13522 14306
rect 13522 14254 13524 14306
rect 13468 14252 13524 14254
rect 18396 17052 18452 17108
rect 18620 17388 18676 17444
rect 18396 15372 18452 15428
rect 19068 18450 19124 18452
rect 19068 18398 19070 18450
rect 19070 18398 19122 18450
rect 19122 18398 19124 18450
rect 19068 18396 19124 18398
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 20860 23772 20916 23828
rect 23548 38220 23604 38276
rect 21532 37436 21588 37492
rect 22764 37490 22820 37492
rect 22764 37438 22766 37490
rect 22766 37438 22818 37490
rect 22818 37438 22820 37490
rect 22764 37436 22820 37438
rect 24220 37436 24276 37492
rect 21084 26908 21140 26964
rect 21644 26962 21700 26964
rect 21644 26910 21646 26962
rect 21646 26910 21698 26962
rect 21698 26910 21700 26962
rect 21644 26908 21700 26910
rect 21308 26796 21364 26852
rect 21308 26402 21364 26404
rect 21308 26350 21310 26402
rect 21310 26350 21362 26402
rect 21362 26350 21364 26402
rect 21308 26348 21364 26350
rect 21084 25228 21140 25284
rect 21644 26402 21700 26404
rect 21644 26350 21646 26402
rect 21646 26350 21698 26402
rect 21698 26350 21700 26402
rect 21644 26348 21700 26350
rect 22316 36706 22372 36708
rect 22316 36654 22318 36706
rect 22318 36654 22370 36706
rect 22370 36654 22372 36706
rect 22316 36652 22372 36654
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 24892 36652 24948 36708
rect 22316 27858 22372 27860
rect 22316 27806 22318 27858
rect 22318 27806 22370 27858
rect 22370 27806 22372 27858
rect 22316 27804 22372 27806
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 22204 27074 22260 27076
rect 22204 27022 22206 27074
rect 22206 27022 22258 27074
rect 22258 27022 22260 27074
rect 22204 27020 22260 27022
rect 23324 27020 23380 27076
rect 22428 26402 22484 26404
rect 22428 26350 22430 26402
rect 22430 26350 22482 26402
rect 22482 26350 22484 26402
rect 22428 26348 22484 26350
rect 21980 25228 22036 25284
rect 21420 23660 21476 23716
rect 19852 20524 19908 20580
rect 20524 20524 20580 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19292 20076 19348 20132
rect 19292 19292 19348 19348
rect 20188 19292 20244 19348
rect 19964 19234 20020 19236
rect 19964 19182 19966 19234
rect 19966 19182 20018 19234
rect 20018 19182 20020 19234
rect 19964 19180 20020 19182
rect 19628 19122 19684 19124
rect 19628 19070 19630 19122
rect 19630 19070 19682 19122
rect 19682 19070 19684 19122
rect 19628 19068 19684 19070
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19292 18060 19348 18116
rect 19180 17500 19236 17556
rect 19852 17778 19908 17780
rect 19852 17726 19854 17778
rect 19854 17726 19906 17778
rect 19906 17726 19908 17778
rect 19852 17724 19908 17726
rect 21420 19852 21476 19908
rect 20748 19234 20804 19236
rect 20748 19182 20750 19234
rect 20750 19182 20802 19234
rect 20802 19182 20804 19234
rect 20748 19180 20804 19182
rect 20860 18284 20916 18340
rect 19964 17612 20020 17668
rect 20076 17836 20132 17892
rect 20300 17388 20356 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20300 17164 20356 17220
rect 20524 17612 20580 17668
rect 19740 17052 19796 17108
rect 19404 16828 19460 16884
rect 20076 17106 20132 17108
rect 20076 17054 20078 17106
rect 20078 17054 20130 17106
rect 20130 17054 20132 17106
rect 20076 17052 20132 17054
rect 21532 19122 21588 19124
rect 21532 19070 21534 19122
rect 21534 19070 21586 19122
rect 21586 19070 21588 19122
rect 21532 19068 21588 19070
rect 21420 18060 21476 18116
rect 21308 17724 21364 17780
rect 21420 17836 21476 17892
rect 18732 15148 18788 15204
rect 19740 16098 19796 16100
rect 19740 16046 19742 16098
rect 19742 16046 19794 16098
rect 19794 16046 19796 16098
rect 19740 16044 19796 16046
rect 20300 16994 20356 16996
rect 20300 16942 20302 16994
rect 20302 16942 20354 16994
rect 20354 16942 20356 16994
rect 20300 16940 20356 16942
rect 20524 16828 20580 16884
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20412 15596 20468 15652
rect 19516 15426 19572 15428
rect 19516 15374 19518 15426
rect 19518 15374 19570 15426
rect 19570 15374 19572 15426
rect 19516 15372 19572 15374
rect 21196 17612 21252 17668
rect 22876 26290 22932 26292
rect 22876 26238 22878 26290
rect 22878 26238 22930 26290
rect 22930 26238 22932 26290
rect 22876 26236 22932 26238
rect 22204 23996 22260 24052
rect 22092 22428 22148 22484
rect 24668 26796 24724 26852
rect 23660 26514 23716 26516
rect 23660 26462 23662 26514
rect 23662 26462 23714 26514
rect 23714 26462 23716 26514
rect 23660 26460 23716 26462
rect 24332 26514 24388 26516
rect 24332 26462 24334 26514
rect 24334 26462 24386 26514
rect 24386 26462 24388 26514
rect 24332 26460 24388 26462
rect 25228 26796 25284 26852
rect 25228 26514 25284 26516
rect 25228 26462 25230 26514
rect 25230 26462 25282 26514
rect 25282 26462 25284 26514
rect 25228 26460 25284 26462
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 26124 36706 26180 36708
rect 26124 36654 26126 36706
rect 26126 36654 26178 36706
rect 26178 36654 26180 36706
rect 26124 36652 26180 36654
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 25676 27074 25732 27076
rect 25676 27022 25678 27074
rect 25678 27022 25730 27074
rect 25730 27022 25732 27074
rect 25676 27020 25732 27022
rect 23436 26290 23492 26292
rect 23436 26238 23438 26290
rect 23438 26238 23490 26290
rect 23490 26238 23492 26290
rect 23436 26236 23492 26238
rect 22428 23154 22484 23156
rect 22428 23102 22430 23154
rect 22430 23102 22482 23154
rect 22482 23102 22484 23154
rect 22428 23100 22484 23102
rect 23212 23100 23268 23156
rect 22316 22540 22372 22596
rect 22764 22428 22820 22484
rect 22652 20802 22708 20804
rect 22652 20750 22654 20802
rect 22654 20750 22706 20802
rect 22706 20750 22708 20802
rect 22652 20748 22708 20750
rect 22540 19010 22596 19012
rect 22540 18958 22542 19010
rect 22542 18958 22594 19010
rect 22594 18958 22596 19010
rect 22540 18956 22596 18958
rect 21980 18396 22036 18452
rect 21756 17948 21812 18004
rect 21420 17164 21476 17220
rect 22204 17500 22260 17556
rect 21756 17164 21812 17220
rect 21532 17052 21588 17108
rect 23324 22370 23380 22372
rect 23324 22318 23326 22370
rect 23326 22318 23378 22370
rect 23378 22318 23380 22370
rect 23324 22316 23380 22318
rect 23324 22092 23380 22148
rect 22876 20524 22932 20580
rect 22652 17724 22708 17780
rect 22316 17164 22372 17220
rect 20860 16044 20916 16100
rect 22316 15484 22372 15540
rect 22428 15596 22484 15652
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 16940 13356 16996 13412
rect 4684 13300 4740 13302
rect 15820 13074 15876 13076
rect 15820 13022 15822 13074
rect 15822 13022 15874 13074
rect 15874 13022 15876 13074
rect 15820 13020 15876 13022
rect 17948 13356 18004 13412
rect 17500 13020 17556 13076
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18620 13356 18676 13412
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20860 3612 20916 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21644 14306 21700 14308
rect 21644 14254 21646 14306
rect 21646 14254 21698 14306
rect 21698 14254 21700 14306
rect 21644 14252 21700 14254
rect 23324 19234 23380 19236
rect 23324 19182 23326 19234
rect 23326 19182 23378 19234
rect 23378 19182 23380 19234
rect 23324 19180 23380 19182
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 25900 23266 25956 23268
rect 25900 23214 25902 23266
rect 25902 23214 25954 23266
rect 25954 23214 25956 23266
rect 25900 23212 25956 23214
rect 25340 23100 25396 23156
rect 24332 23042 24388 23044
rect 24332 22990 24334 23042
rect 24334 22990 24386 23042
rect 24386 22990 24388 23042
rect 24332 22988 24388 22990
rect 24108 22428 24164 22484
rect 24444 22876 24500 22932
rect 23884 22204 23940 22260
rect 23772 22092 23828 22148
rect 25340 22930 25396 22932
rect 25340 22878 25342 22930
rect 25342 22878 25394 22930
rect 25394 22878 25396 22930
rect 25340 22876 25396 22878
rect 25228 22316 25284 22372
rect 26236 23100 26292 23156
rect 25900 22988 25956 23044
rect 26236 22482 26292 22484
rect 26236 22430 26238 22482
rect 26238 22430 26290 22482
rect 26290 22430 26292 22482
rect 26236 22428 26292 22430
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 40012 23548 40068 23604
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 37884 22428 37940 22484
rect 26572 22316 26628 22372
rect 25452 22092 25508 22148
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 23548 18844 23604 18900
rect 23548 18508 23604 18564
rect 23212 18172 23268 18228
rect 23212 17612 23268 17668
rect 23436 17836 23492 17892
rect 23660 18284 23716 18340
rect 24108 19964 24164 20020
rect 25676 20018 25732 20020
rect 25676 19966 25678 20018
rect 25678 19966 25730 20018
rect 25730 19966 25732 20018
rect 25676 19964 25732 19966
rect 24332 18844 24388 18900
rect 24556 18674 24612 18676
rect 24556 18622 24558 18674
rect 24558 18622 24610 18674
rect 24610 18622 24612 18674
rect 24556 18620 24612 18622
rect 24108 18562 24164 18564
rect 24108 18510 24110 18562
rect 24110 18510 24162 18562
rect 24162 18510 24164 18562
rect 24108 18508 24164 18510
rect 24668 18508 24724 18564
rect 23884 18172 23940 18228
rect 24668 18172 24724 18228
rect 23548 17612 23604 17668
rect 23436 17554 23492 17556
rect 23436 17502 23438 17554
rect 23438 17502 23490 17554
rect 23490 17502 23492 17554
rect 23436 17500 23492 17502
rect 25004 18508 25060 18564
rect 29036 20018 29092 20020
rect 29036 19966 29038 20018
rect 29038 19966 29090 20018
rect 29090 19966 29092 20018
rect 29036 19964 29092 19966
rect 26012 18956 26068 19012
rect 27916 19852 27972 19908
rect 29484 19906 29540 19908
rect 29484 19854 29486 19906
rect 29486 19854 29538 19906
rect 29538 19854 29540 19906
rect 29484 19852 29540 19854
rect 26908 19180 26964 19236
rect 27356 19180 27412 19236
rect 26236 19068 26292 19124
rect 27132 18620 27188 18676
rect 27020 18562 27076 18564
rect 27020 18510 27022 18562
rect 27022 18510 27074 18562
rect 27074 18510 27076 18562
rect 27020 18508 27076 18510
rect 26796 18450 26852 18452
rect 26796 18398 26798 18450
rect 26798 18398 26850 18450
rect 26850 18398 26852 18450
rect 26796 18396 26852 18398
rect 26124 18284 26180 18340
rect 26460 18284 26516 18340
rect 25788 18172 25844 18228
rect 27132 18338 27188 18340
rect 27132 18286 27134 18338
rect 27134 18286 27186 18338
rect 27186 18286 27188 18338
rect 27132 18284 27188 18286
rect 27020 18172 27076 18228
rect 24108 17554 24164 17556
rect 24108 17502 24110 17554
rect 24110 17502 24162 17554
rect 24162 17502 24164 17554
rect 24108 17500 24164 17502
rect 23324 15484 23380 15540
rect 24892 17554 24948 17556
rect 24892 17502 24894 17554
rect 24894 17502 24946 17554
rect 24946 17502 24948 17554
rect 24892 17500 24948 17502
rect 23548 15314 23604 15316
rect 23548 15262 23550 15314
rect 23550 15262 23602 15314
rect 23602 15262 23604 15314
rect 23548 15260 23604 15262
rect 22316 15036 22372 15092
rect 22540 15090 22596 15092
rect 22540 15038 22542 15090
rect 22542 15038 22594 15090
rect 22594 15038 22596 15090
rect 22540 15036 22596 15038
rect 22204 14252 22260 14308
rect 22652 14306 22708 14308
rect 22652 14254 22654 14306
rect 22654 14254 22706 14306
rect 22706 14254 22708 14306
rect 22652 14252 22708 14254
rect 28924 19068 28980 19124
rect 27356 18172 27412 18228
rect 26684 16994 26740 16996
rect 26684 16942 26686 16994
rect 26686 16942 26738 16994
rect 26738 16942 26740 16994
rect 26684 16940 26740 16942
rect 27804 17612 27860 17668
rect 28588 17612 28644 17668
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 20860 40068 20916
rect 37884 19964 37940 20020
rect 40012 19516 40068 19572
rect 37660 19180 37716 19236
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 27244 16828 27300 16884
rect 28588 16828 28644 16884
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 17500 40068 17556
rect 37660 16882 37716 16884
rect 37660 16830 37662 16882
rect 37662 16830 37714 16882
rect 37714 16830 37716 16882
rect 37660 16828 37716 16830
rect 40012 16828 40068 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 24444 14700 24500 14756
rect 25564 14700 25620 14756
rect 24556 14588 24612 14644
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 25676 14588 25732 14644
rect 26348 14588 26404 14644
rect 26908 14642 26964 14644
rect 26908 14590 26910 14642
rect 26910 14590 26962 14642
rect 26962 14590 26964 14642
rect 26908 14588 26964 14590
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 15362 38220 15372 38276
rect 15428 38220 16156 38276
rect 16212 38220 16222 38276
rect 23538 38220 23548 38276
rect 23604 38220 25564 38276
rect 25620 38220 25630 38276
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 21522 37436 21532 37492
rect 21588 37436 22764 37492
rect 22820 37436 22830 37492
rect 24210 37436 24220 37492
rect 24276 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 16818 36652 16828 36708
rect 16884 36652 18060 36708
rect 18116 36652 18126 36708
rect 20850 36652 20860 36708
rect 20916 36652 22316 36708
rect 22372 36652 22382 36708
rect 24882 36652 24892 36708
rect 24948 36652 26124 36708
rect 26180 36652 26190 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 13794 28028 13804 28084
rect 13860 28028 14812 28084
rect 14868 28028 14878 28084
rect 15026 27804 15036 27860
rect 15092 27804 16044 27860
rect 16100 27804 16110 27860
rect 18946 27804 18956 27860
rect 19012 27804 22316 27860
rect 22372 27804 22382 27860
rect 15026 27580 15036 27636
rect 15092 27580 16044 27636
rect 16100 27580 16110 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 16258 27132 16268 27188
rect 16324 27132 17164 27188
rect 17220 27132 17230 27188
rect 19506 27132 19516 27188
rect 19572 27132 20524 27188
rect 20580 27132 20590 27188
rect 4274 27020 4284 27076
rect 4340 27020 11228 27076
rect 11284 27020 14140 27076
rect 14196 27020 14206 27076
rect 22194 27020 22204 27076
rect 22260 27020 23324 27076
rect 23380 27020 25676 27076
rect 25732 27020 25742 27076
rect 0 26964 800 26992
rect 0 26908 4172 26964
rect 4228 26908 4238 26964
rect 14242 26908 14252 26964
rect 14308 26908 14318 26964
rect 21074 26908 21084 26964
rect 21140 26908 21644 26964
rect 21700 26908 21710 26964
rect 0 26880 800 26908
rect 14252 26852 14308 26908
rect 13122 26796 13132 26852
rect 13188 26796 14308 26852
rect 15586 26796 15596 26852
rect 15652 26796 16604 26852
rect 16660 26796 16670 26852
rect 19618 26796 19628 26852
rect 19684 26796 20748 26852
rect 20804 26796 20814 26852
rect 21298 26796 21308 26852
rect 21364 26796 21374 26852
rect 24658 26796 24668 26852
rect 24724 26796 25228 26852
rect 25284 26796 25294 26852
rect 16146 26684 16156 26740
rect 16212 26684 18844 26740
rect 18900 26684 18910 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 16706 26460 16716 26516
rect 16772 26460 18508 26516
rect 18564 26460 18574 26516
rect 21308 26404 21364 26796
rect 23650 26460 23660 26516
rect 23716 26460 24332 26516
rect 24388 26460 25228 26516
rect 25284 26460 25294 26516
rect 17612 26348 19964 26404
rect 20020 26348 21308 26404
rect 21364 26348 21374 26404
rect 21634 26348 21644 26404
rect 21700 26348 22428 26404
rect 22484 26348 22494 26404
rect 0 26292 800 26320
rect 17612 26292 17668 26348
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 16818 26236 16828 26292
rect 16884 26236 17612 26292
rect 17668 26236 17678 26292
rect 18834 26236 18844 26292
rect 18900 26236 19852 26292
rect 19908 26236 20412 26292
rect 20468 26236 20478 26292
rect 0 26208 800 26236
rect 21644 26180 21700 26348
rect 22866 26236 22876 26292
rect 22932 26236 23436 26292
rect 23492 26236 23502 26292
rect 16594 26124 16604 26180
rect 16660 26124 21700 26180
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 13346 25676 13356 25732
rect 13412 25676 14812 25732
rect 14868 25676 14878 25732
rect 15138 25676 15148 25732
rect 15204 25676 15214 25732
rect 15148 25620 15204 25676
rect 15148 25564 15372 25620
rect 15428 25564 15438 25620
rect 15138 25452 15148 25508
rect 15204 25452 16604 25508
rect 16660 25452 16670 25508
rect 14130 25340 14140 25396
rect 14196 25340 14812 25396
rect 14868 25340 16492 25396
rect 16548 25340 16558 25396
rect 13122 25228 13132 25284
rect 13188 25228 14364 25284
rect 14420 25228 16268 25284
rect 16324 25228 17500 25284
rect 17556 25228 17566 25284
rect 19058 25228 19068 25284
rect 19124 25228 20636 25284
rect 20692 25228 21084 25284
rect 21140 25228 21980 25284
rect 22036 25228 22046 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 14914 23996 14924 24052
rect 14980 23996 15932 24052
rect 15988 23996 22204 24052
rect 22260 23996 22270 24052
rect 4274 23884 4284 23940
rect 4340 23884 8428 23940
rect 16706 23884 16716 23940
rect 16772 23884 17836 23940
rect 17892 23884 17902 23940
rect 8372 23828 8428 23884
rect 8372 23772 11004 23828
rect 11060 23772 14364 23828
rect 14420 23772 14430 23828
rect 15698 23772 15708 23828
rect 15764 23772 17276 23828
rect 17332 23772 19068 23828
rect 19124 23772 19134 23828
rect 19394 23772 19404 23828
rect 19460 23772 20636 23828
rect 20692 23772 20860 23828
rect 20916 23772 20926 23828
rect 14242 23660 14252 23716
rect 14308 23660 15596 23716
rect 15652 23660 15662 23716
rect 19842 23660 19852 23716
rect 19908 23660 21420 23716
rect 21476 23660 21486 23716
rect 0 23604 800 23632
rect 41200 23604 42000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 17602 23436 17612 23492
rect 17668 23436 19628 23492
rect 19684 23436 19694 23492
rect 25890 23212 25900 23268
rect 25956 23212 31948 23268
rect 31892 23156 31948 23212
rect 4274 23100 4284 23156
rect 4340 23100 13692 23156
rect 13748 23100 15708 23156
rect 15764 23100 15774 23156
rect 18946 23100 18956 23156
rect 19012 23100 22428 23156
rect 22484 23100 23212 23156
rect 23268 23100 23278 23156
rect 25330 23100 25340 23156
rect 25396 23100 26236 23156
rect 26292 23100 26302 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 13570 22988 13580 23044
rect 13636 22988 13916 23044
rect 13972 22988 16492 23044
rect 16548 22988 16940 23044
rect 16996 22988 17500 23044
rect 17556 22988 17566 23044
rect 24322 22988 24332 23044
rect 24388 22988 25900 23044
rect 25956 22988 25966 23044
rect 0 22932 800 22960
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 24434 22876 24444 22932
rect 24500 22876 25340 22932
rect 25396 22876 25406 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 13122 22540 13132 22596
rect 13188 22540 13916 22596
rect 13972 22540 13982 22596
rect 17714 22540 17724 22596
rect 17780 22540 18508 22596
rect 18564 22540 22316 22596
rect 22372 22540 22382 22596
rect 1922 22428 1932 22484
rect 1988 22428 1998 22484
rect 8372 22428 9996 22484
rect 10052 22428 14588 22484
rect 14644 22428 14654 22484
rect 15586 22428 15596 22484
rect 15652 22428 17612 22484
rect 17668 22428 17678 22484
rect 22082 22428 22092 22484
rect 22148 22428 22764 22484
rect 22820 22428 24108 22484
rect 24164 22428 24174 22484
rect 26226 22428 26236 22484
rect 26292 22428 37884 22484
rect 37940 22428 37950 22484
rect 0 22260 800 22288
rect 1932 22260 1988 22428
rect 8372 22372 8428 22428
rect 4274 22316 4284 22372
rect 4340 22316 8428 22372
rect 12898 22316 12908 22372
rect 12964 22316 13580 22372
rect 13636 22316 13646 22372
rect 14466 22316 14476 22372
rect 14532 22316 15036 22372
rect 15092 22316 16212 22372
rect 16594 22316 16604 22372
rect 16660 22316 17388 22372
rect 17444 22316 17454 22372
rect 23314 22316 23324 22372
rect 23380 22316 25228 22372
rect 25284 22316 26572 22372
rect 26628 22316 26638 22372
rect 16156 22260 16212 22316
rect 0 22204 1988 22260
rect 16146 22204 16156 22260
rect 16212 22204 16222 22260
rect 19506 22204 19516 22260
rect 19572 22204 20860 22260
rect 20916 22204 23884 22260
rect 23940 22204 23950 22260
rect 0 22176 800 22204
rect 15810 22092 15820 22148
rect 15876 22092 16492 22148
rect 16548 22092 16558 22148
rect 23314 22092 23324 22148
rect 23380 22092 23772 22148
rect 23828 22092 25452 22148
rect 25508 22092 25518 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 12114 21756 12124 21812
rect 12180 21756 14700 21812
rect 14756 21756 14766 21812
rect 15810 21756 15820 21812
rect 15876 21756 18396 21812
rect 18452 21756 19292 21812
rect 19348 21756 19358 21812
rect 16818 21644 16828 21700
rect 16884 21644 19404 21700
rect 19460 21644 19964 21700
rect 20020 21644 20030 21700
rect 15474 21532 15484 21588
rect 15540 21532 19852 21588
rect 19908 21532 19918 21588
rect 4162 21420 4172 21476
rect 4228 21420 18060 21476
rect 18116 21420 18956 21476
rect 19012 21420 19022 21476
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 15026 21084 15036 21140
rect 15092 21084 15820 21140
rect 15876 21084 15886 21140
rect 41200 20916 42000 20944
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 20066 20748 20076 20804
rect 20132 20748 22652 20804
rect 22708 20748 22718 20804
rect 19842 20524 19852 20580
rect 19908 20524 20524 20580
rect 20580 20524 22876 20580
rect 22932 20524 22942 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 14690 20076 14700 20132
rect 14756 20076 15484 20132
rect 15540 20076 15550 20132
rect 17826 20076 17836 20132
rect 17892 20076 18508 20132
rect 18564 20076 19292 20132
rect 19348 20076 19358 20132
rect 13906 19964 13916 20020
rect 13972 19964 16156 20020
rect 16212 19964 18284 20020
rect 18340 19964 18350 20020
rect 24098 19964 24108 20020
rect 24164 19964 25676 20020
rect 25732 19964 26908 20020
rect 29026 19964 29036 20020
rect 29092 19964 37884 20020
rect 37940 19964 37950 20020
rect 26852 19908 26908 19964
rect 17938 19852 17948 19908
rect 18004 19852 18844 19908
rect 18900 19852 21420 19908
rect 21476 19852 21486 19908
rect 26852 19852 27916 19908
rect 27972 19852 29484 19908
rect 29540 19852 29550 19908
rect 18172 19796 18228 19852
rect 18162 19740 18172 19796
rect 18228 19740 18238 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 15250 19292 15260 19348
rect 15316 19292 16604 19348
rect 16660 19292 16670 19348
rect 19282 19292 19292 19348
rect 19348 19292 20188 19348
rect 20244 19292 20254 19348
rect 4274 19180 4284 19236
rect 4340 19180 8428 19236
rect 16706 19180 16716 19236
rect 16772 19180 18172 19236
rect 18228 19180 18238 19236
rect 18722 19180 18732 19236
rect 18788 19180 19068 19236
rect 19124 19180 19964 19236
rect 20020 19180 20030 19236
rect 20738 19180 20748 19236
rect 20804 19180 23324 19236
rect 23380 19180 23390 19236
rect 26898 19180 26908 19236
rect 26964 19180 27356 19236
rect 27412 19180 37660 19236
rect 37716 19180 37726 19236
rect 8372 19012 8428 19180
rect 11778 19068 11788 19124
rect 11844 19068 14924 19124
rect 14980 19068 14990 19124
rect 16930 19068 16940 19124
rect 16996 19068 17276 19124
rect 17332 19068 17342 19124
rect 17602 19068 17612 19124
rect 17668 19068 19460 19124
rect 19618 19068 19628 19124
rect 19684 19068 21532 19124
rect 21588 19068 21598 19124
rect 26226 19068 26236 19124
rect 26292 19068 28924 19124
rect 28980 19068 28990 19124
rect 19404 19012 19460 19068
rect 8372 18956 9996 19012
rect 10052 18956 14252 19012
rect 14308 18956 14318 19012
rect 15362 18956 15372 19012
rect 15428 18956 17500 19012
rect 17556 18956 17566 19012
rect 19404 18956 22372 19012
rect 22530 18956 22540 19012
rect 22596 18956 26012 19012
rect 26068 18956 26078 19012
rect 0 18900 800 18928
rect 22316 18900 22372 18956
rect 0 18844 1932 18900
rect 1988 18844 1998 18900
rect 22316 18844 23548 18900
rect 23604 18844 24332 18900
rect 24388 18844 24398 18900
rect 0 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 14018 18620 14028 18676
rect 14084 18620 17948 18676
rect 18004 18620 24388 18676
rect 24546 18620 24556 18676
rect 24612 18620 27132 18676
rect 27188 18620 27198 18676
rect 24332 18564 24388 18620
rect 17266 18508 17276 18564
rect 17332 18508 23548 18564
rect 23604 18508 24108 18564
rect 24164 18508 24174 18564
rect 24332 18508 24668 18564
rect 24724 18508 24734 18564
rect 24994 18508 25004 18564
rect 25060 18508 27020 18564
rect 27076 18508 27086 18564
rect 11106 18396 11116 18452
rect 11172 18396 12796 18452
rect 12852 18396 12862 18452
rect 15922 18396 15932 18452
rect 15988 18396 16156 18452
rect 16212 18396 16222 18452
rect 18162 18396 18172 18452
rect 18228 18396 19068 18452
rect 19124 18396 19134 18452
rect 21970 18396 21980 18452
rect 22036 18396 26796 18452
rect 26852 18396 26862 18452
rect 15474 18284 15484 18340
rect 15540 18284 16380 18340
rect 16436 18284 16446 18340
rect 17602 18284 17612 18340
rect 17668 18284 18732 18340
rect 18788 18284 18798 18340
rect 20822 18284 20860 18340
rect 20916 18284 20926 18340
rect 23650 18284 23660 18340
rect 23716 18284 26124 18340
rect 26180 18284 26190 18340
rect 26450 18284 26460 18340
rect 26516 18284 27132 18340
rect 27188 18284 27198 18340
rect 26124 18228 26180 18284
rect 12114 18172 12124 18228
rect 12180 18172 14700 18228
rect 14756 18172 14766 18228
rect 16482 18172 16492 18228
rect 16548 18172 18284 18228
rect 18340 18172 18350 18228
rect 18498 18172 18508 18228
rect 18564 18172 23212 18228
rect 23268 18172 23884 18228
rect 23940 18172 23950 18228
rect 24658 18172 24668 18228
rect 24724 18172 25788 18228
rect 25844 18172 25854 18228
rect 26124 18172 27020 18228
rect 27076 18172 27356 18228
rect 27412 18172 27422 18228
rect 16370 18060 16380 18116
rect 16436 18060 17612 18116
rect 17668 18060 17678 18116
rect 17938 18060 17948 18116
rect 18004 18060 19292 18116
rect 19348 18060 21420 18116
rect 21476 18060 21486 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 16706 17948 16716 18004
rect 16772 17948 21756 18004
rect 21812 17948 21822 18004
rect 17154 17836 17164 17892
rect 17220 17836 18396 17892
rect 18452 17836 18462 17892
rect 20066 17836 20076 17892
rect 20132 17836 21420 17892
rect 21476 17836 23436 17892
rect 23492 17836 23502 17892
rect 16258 17724 16268 17780
rect 16324 17724 19852 17780
rect 19908 17724 21308 17780
rect 21364 17724 21374 17780
rect 22642 17724 22652 17780
rect 22708 17724 24164 17780
rect 12786 17612 12796 17668
rect 12852 17612 13580 17668
rect 13636 17612 14140 17668
rect 14196 17612 14206 17668
rect 16482 17612 16492 17668
rect 16548 17612 17164 17668
rect 17220 17612 17230 17668
rect 17378 17612 17388 17668
rect 17444 17612 18060 17668
rect 18116 17612 19964 17668
rect 20020 17612 20524 17668
rect 20580 17612 21196 17668
rect 21252 17612 21262 17668
rect 23202 17612 23212 17668
rect 23268 17612 23548 17668
rect 23604 17612 23614 17668
rect 24108 17556 24164 17724
rect 27794 17612 27804 17668
rect 27860 17612 28588 17668
rect 28644 17612 37660 17668
rect 37716 17612 37726 17668
rect 41200 17556 42000 17584
rect 15810 17500 15820 17556
rect 15876 17500 17500 17556
rect 17556 17500 17566 17556
rect 18274 17500 18284 17556
rect 18340 17500 19180 17556
rect 19236 17500 19246 17556
rect 22194 17500 22204 17556
rect 22260 17500 23436 17556
rect 23492 17500 23502 17556
rect 24098 17500 24108 17556
rect 24164 17500 24892 17556
rect 24948 17500 24958 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 14690 17388 14700 17444
rect 14756 17388 15372 17444
rect 15428 17388 16492 17444
rect 16548 17388 16558 17444
rect 18610 17388 18620 17444
rect 18676 17388 20300 17444
rect 20356 17388 20366 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 20290 17164 20300 17220
rect 20356 17164 21420 17220
rect 21476 17164 21756 17220
rect 21812 17164 22316 17220
rect 22372 17164 22382 17220
rect 17602 17052 17612 17108
rect 17668 17052 18396 17108
rect 18452 17052 19740 17108
rect 19796 17052 19806 17108
rect 20066 17052 20076 17108
rect 20132 17052 21532 17108
rect 21588 17052 21598 17108
rect 20290 16940 20300 16996
rect 20356 16940 26684 16996
rect 26740 16940 26750 16996
rect 41200 16884 42000 16912
rect 12786 16828 12796 16884
rect 12852 16828 14028 16884
rect 14084 16828 14094 16884
rect 19394 16828 19404 16884
rect 19460 16828 20524 16884
rect 20580 16828 20590 16884
rect 27234 16828 27244 16884
rect 27300 16828 28588 16884
rect 28644 16828 37660 16884
rect 37716 16828 37726 16884
rect 40002 16828 40012 16884
rect 40068 16828 42000 16884
rect 41200 16800 42000 16828
rect 15586 16716 15596 16772
rect 15652 16716 17500 16772
rect 17556 16716 17566 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16212 800 16240
rect 0 16156 1932 16212
rect 1988 16156 1998 16212
rect 0 16128 800 16156
rect 19730 16044 19740 16100
rect 19796 16044 20860 16100
rect 20916 16044 20926 16100
rect 4274 15708 4284 15764
rect 4340 15708 10668 15764
rect 10724 15708 13692 15764
rect 13748 15708 13758 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 20402 15596 20412 15652
rect 20468 15596 22428 15652
rect 22484 15596 22494 15652
rect 0 15540 800 15568
rect 0 15484 2044 15540
rect 2100 15484 2110 15540
rect 22306 15484 22316 15540
rect 22372 15484 22540 15540
rect 22596 15484 23324 15540
rect 23380 15484 23390 15540
rect 0 15456 800 15484
rect 4274 15372 4284 15428
rect 4340 15372 13468 15428
rect 13524 15372 13534 15428
rect 18386 15372 18396 15428
rect 18452 15372 19516 15428
rect 19572 15372 19582 15428
rect 13570 15260 13580 15316
rect 13636 15260 13916 15316
rect 13972 15260 16940 15316
rect 16996 15260 17500 15316
rect 17556 15260 17566 15316
rect 22316 15260 23548 15316
rect 23604 15260 23614 15316
rect 16818 15148 16828 15204
rect 16884 15148 18732 15204
rect 18788 15148 18798 15204
rect 22316 15092 22372 15260
rect 22530 15148 22540 15204
rect 22596 15148 22606 15204
rect 22540 15092 22596 15148
rect 1922 15036 1932 15092
rect 1988 15036 1998 15092
rect 22306 15036 22316 15092
rect 22372 15036 22382 15092
rect 22530 15036 22540 15092
rect 22596 15036 22606 15092
rect 0 14868 800 14896
rect 1932 14868 1988 15036
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 0 14812 1988 14868
rect 0 14784 800 14812
rect 24434 14700 24444 14756
rect 24500 14700 25564 14756
rect 25620 14700 25630 14756
rect 24546 14588 24556 14644
rect 24612 14588 25676 14644
rect 25732 14588 26348 14644
rect 26404 14588 26908 14644
rect 26964 14588 26974 14644
rect 4050 14252 4060 14308
rect 4116 14252 13468 14308
rect 13524 14252 13534 14308
rect 21634 14252 21644 14308
rect 21700 14252 22204 14308
rect 22260 14252 22652 14308
rect 22708 14252 22718 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 16930 13356 16940 13412
rect 16996 13356 17948 13412
rect 18004 13356 18620 13412
rect 18676 13356 18686 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 15810 13020 15820 13076
rect 15876 13020 17500 13076
rect 17556 13020 17566 13076
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 20860 22204 20916 22260
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 20860 18284 20916 18340
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 22540 15484 22596 15540
rect 22540 15148 22596 15204
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 20860 22260 20916 22270
rect 20860 18340 20916 22204
rect 20860 18274 20916 18284
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 22540 15540 22596 15550
rect 22540 15204 22596 15484
rect 22540 15138 22596 15148
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _099_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _102_
timestamp 1698175906
transform -1 0 22848 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21840 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21728 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform 1 0 16016 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_
timestamp 1698175906
transform -1 0 18144 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _107_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _108_
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 19152 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform -1 0 20384 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22512 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _114_
timestamp 1698175906
transform -1 0 22512 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23072 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _116_
timestamp 1698175906
transform 1 0 20608 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _118_
timestamp 1698175906
transform 1 0 18480 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 21728 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 20384 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform -1 0 20832 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _123_
timestamp 1698175906
transform 1 0 18144 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _124_
timestamp 1698175906
transform 1 0 19376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _125_
timestamp 1698175906
transform -1 0 22736 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20832 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _127_
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform -1 0 18928 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20160 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23072 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1698175906
transform 1 0 23968 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 23744 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform 1 0 23296 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1698175906
transform -1 0 17136 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 15792 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15680 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _138_
timestamp 1698175906
transform -1 0 16016 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _139_
timestamp 1698175906
transform -1 0 16912 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _141_
timestamp 1698175906
transform -1 0 15792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 19824 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _143_
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform 1 0 23184 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 27552 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 26992 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform 1 0 18928 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _149_
timestamp 1698175906
transform -1 0 20160 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform -1 0 16016 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19264 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _152_
timestamp 1698175906
transform -1 0 20160 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform -1 0 18144 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 27664 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _155_
timestamp 1698175906
transform 1 0 23968 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _156_
timestamp 1698175906
transform 1 0 21168 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22512 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 23968 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _159_
timestamp 1698175906
transform 1 0 22064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform 1 0 25648 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24528 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 25648 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _163_
timestamp 1698175906
transform -1 0 24640 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _165_
timestamp 1698175906
transform -1 0 17024 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _166_
timestamp 1698175906
transform -1 0 16352 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _167_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15904 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _168_
timestamp 1698175906
transform -1 0 29232 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _169_
timestamp 1698175906
transform 1 0 22176 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1698175906
transform -1 0 18480 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _171_
timestamp 1698175906
transform 1 0 25648 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _172_
timestamp 1698175906
transform 1 0 14000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _173_
timestamp 1698175906
transform -1 0 15344 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _174_
timestamp 1698175906
transform 1 0 13776 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _175_
timestamp 1698175906
transform -1 0 17808 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _176_
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _177_
timestamp 1698175906
transform 1 0 14448 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform 1 0 14000 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _179_
timestamp 1698175906
transform 1 0 14560 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1698175906
transform 1 0 17360 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _181_
timestamp 1698175906
transform -1 0 18592 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _182_
timestamp 1698175906
transform -1 0 18480 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _183_
timestamp 1698175906
transform -1 0 16912 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _184_
timestamp 1698175906
transform 1 0 15792 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _185_
timestamp 1698175906
transform -1 0 16016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _186_
timestamp 1698175906
transform -1 0 15792 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform 1 0 15456 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1698175906
transform -1 0 17920 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _189_
timestamp 1698175906
transform 1 0 16016 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform -1 0 14672 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16352 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 14448 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _193_
timestamp 1698175906
transform -1 0 28000 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _194_
timestamp 1698175906
transform 1 0 24304 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _195_
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _197_
timestamp 1698175906
transform 1 0 26656 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 17472 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 17808 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform -1 0 24304 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform -1 0 26656 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 10864 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 13776 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 25536 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _206_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18704 0 -1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 23856 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _208_
timestamp 1698175906
transform 1 0 21952 0 1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 23072 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 23184 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform -1 0 13104 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 25536 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 13776 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform -1 0 13104 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform -1 0 14336 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform -1 0 18928 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 14112 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 12880 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform -1 0 16800 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform -1 0 14112 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 25536 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _222_
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _223_
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _224_
timestamp 1698175906
transform -1 0 14000 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _225_
timestamp 1698175906
transform 1 0 24192 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _226_
timestamp 1698175906
transform -1 0 14000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _227_
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A1
timestamp 1698175906
transform 1 0 21952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__A1
timestamp 1698175906
transform 1 0 17248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__A1
timestamp 1698175906
transform 1 0 24080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform -1 0 22400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 26880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 14112 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 29232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 22400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 27888 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 25648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 26544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 26656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 29456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform -1 0 14560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 19152 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 16240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 14336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18816 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20832 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22512 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_123
timestamp 1698175906
transform 1 0 15120 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_127
timestamp 1698175906
transform 1 0 15568 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_157
timestamp 1698175906
transform 1 0 18928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_161 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_169
timestamp 1698175906
transform 1 0 20272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698175906
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_205
timestamp 1698175906
transform 1 0 24304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_113
timestamp 1698175906
transform 1 0 14000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_117
timestamp 1698175906
transform 1 0 14448 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_133
timestamp 1698175906
transform 1 0 16240 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_141
timestamp 1698175906
transform 1 0 17136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_153
timestamp 1698175906
transform 1 0 18480 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_169
timestamp 1698175906
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_226
timestamp 1698175906
transform 1 0 26656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_230
timestamp 1698175906
transform 1 0 27104 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_238
timestamp 1698175906
transform 1 0 28000 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_28
timestamp 1698175906
transform 1 0 4480 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_60
timestamp 1698175906
transform 1 0 8064 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698175906
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_80
timestamp 1698175906
transform 1 0 10304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_154
timestamp 1698175906
transform 1 0 18592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_158
timestamp 1698175906
transform 1 0 19040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_160
timestamp 1698175906
transform 1 0 19264 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_174
timestamp 1698175906
transform 1 0 20832 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_182
timestamp 1698175906
transform 1 0 21728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_184
timestamp 1698175906
transform 1 0 21952 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_191
timestamp 1698175906
transform 1 0 22736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_193
timestamp 1698175906
transform 1 0 22960 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 4480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_117
timestamp 1698175906
transform 1 0 14448 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_121
timestamp 1698175906
transform 1 0 14896 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_129
timestamp 1698175906
transform 1 0 15792 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_145
timestamp 1698175906
transform 1 0 17584 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_149
timestamp 1698175906
transform 1 0 18032 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_195
timestamp 1698175906
transform 1 0 23184 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_199
timestamp 1698175906
transform 1 0 23632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_201
timestamp 1698175906
transform 1 0 23856 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_208
timestamp 1698175906
transform 1 0 24640 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_251
timestamp 1698175906
transform 1 0 29456 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 4480 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1698175906
transform 1 0 13440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698175906
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_121
timestamp 1698175906
transform 1 0 14896 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_148
timestamp 1698175906
transform 1 0 17920 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_164
timestamp 1698175906
transform 1 0 19712 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_182
timestamp 1698175906
transform 1 0 21728 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_192
timestamp 1698175906
transform 1 0 22848 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698175906
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_238
timestamp 1698175906
transform 1 0 28000 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_270
timestamp 1698175906
transform 1 0 31584 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 37408 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_69
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_73
timestamp 1698175906
transform 1 0 9520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_75
timestamp 1698175906
transform 1 0 9744 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_113
timestamp 1698175906
transform 1 0 14000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_116
timestamp 1698175906
transform 1 0 14336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_118
timestamp 1698175906
transform 1 0 14560 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_139
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_143
timestamp 1698175906
transform 1 0 17360 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_154
timestamp 1698175906
transform 1 0 18592 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_183
timestamp 1698175906
transform 1 0 21840 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_191
timestamp 1698175906
transform 1 0 22736 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_195
timestamp 1698175906
transform 1 0 23184 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_201
timestamp 1698175906
transform 1 0 23856 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_212
timestamp 1698175906
transform 1 0 25088 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_251
timestamp 1698175906
transform 1 0 29456 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_84
timestamp 1698175906
transform 1 0 10752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_114
timestamp 1698175906
transform 1 0 14112 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_116
timestamp 1698175906
transform 1 0 14336 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_128
timestamp 1698175906
transform 1 0 15680 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_200
timestamp 1698175906
transform 1 0 23744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_216
timestamp 1698175906
transform 1 0 25536 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_235
timestamp 1698175906
transform 1 0 27664 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_267
timestamp 1698175906
transform 1 0 31248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_275
timestamp 1698175906
transform 1 0 32144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_111
timestamp 1698175906
transform 1 0 13776 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_134
timestamp 1698175906
transform 1 0 16352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_183
timestamp 1698175906
transform 1 0 21840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698175906
transform 1 0 22064 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_194
timestamp 1698175906
transform 1 0 23072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_235
timestamp 1698175906
transform 1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_239
timestamp 1698175906
transform 1 0 28112 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_120
timestamp 1698175906
transform 1 0 14784 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_124
timestamp 1698175906
transform 1 0 15232 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 17472 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698175906
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_249
timestamp 1698175906
transform 1 0 29232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_253
timestamp 1698175906
transform 1 0 29680 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_269
timestamp 1698175906
transform 1 0 31472 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698175906
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_123
timestamp 1698175906
transform 1 0 15120 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_182
timestamp 1698175906
transform 1 0 21728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_186
timestamp 1698175906
transform 1 0 22176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_188
timestamp 1698175906
transform 1 0 22400 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_239
timestamp 1698175906
transform 1 0 28112 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_104
timestamp 1698175906
transform 1 0 12992 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_112
timestamp 1698175906
transform 1 0 13888 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_116
timestamp 1698175906
transform 1 0 14336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_118
timestamp 1698175906
transform 1 0 14560 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_130
timestamp 1698175906
transform 1 0 15904 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_138
timestamp 1698175906
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_146
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_148
timestamp 1698175906
transform 1 0 17920 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_168
timestamp 1698175906
transform 1 0 20160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_189
timestamp 1698175906
transform 1 0 22512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698175906
transform 1 0 9744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_121
timestamp 1698175906
transform 1 0 14896 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_125
timestamp 1698175906
transform 1 0 15344 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_148
timestamp 1698175906
transform 1 0 17920 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_156
timestamp 1698175906
transform 1 0 18816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_158
timestamp 1698175906
transform 1 0 19040 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698175906
transform 1 0 20160 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_183
timestamp 1698175906
transform 1 0 21840 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_191
timestamp 1698175906
transform 1 0 22736 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_224
timestamp 1698175906
transform 1 0 26432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_228
timestamp 1698175906
transform 1 0 26880 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_108
timestamp 1698175906
transform 1 0 13440 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_146
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_154
timestamp 1698175906
transform 1 0 18592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_186
timestamp 1698175906
transform 1 0 22176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_190
timestamp 1698175906
transform 1 0 22624 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_194
timestamp 1698175906
transform 1 0 23072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_222
timestamp 1698175906
transform 1 0 26208 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_254
timestamp 1698175906
transform 1 0 29792 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_270
timestamp 1698175906
transform 1 0 31584 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698175906
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_111
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_113
timestamp 1698175906
transform 1 0 14000 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_119
timestamp 1698175906
transform 1 0 14672 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_123
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698175906
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_144
timestamp 1698175906
transform 1 0 17472 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_167
timestamp 1698175906
transform 1 0 20048 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_183
timestamp 1698175906
transform 1 0 21840 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_191
timestamp 1698175906
transform 1 0 22736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_193
timestamp 1698175906
transform 1 0 22960 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_223
timestamp 1698175906
transform 1 0 26320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_227
timestamp 1698175906
transform 1 0 26768 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_84
timestamp 1698175906
transform 1 0 10752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_114
timestamp 1698175906
transform 1 0 14112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_118
timestamp 1698175906
transform 1 0 14560 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_134
timestamp 1698175906
transform 1 0 16352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_150
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_166
timestamp 1698175906
transform 1 0 19936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_170
timestamp 1698175906
transform 1 0 20384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_178
timestamp 1698175906
transform 1 0 21280 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_111
timestamp 1698175906
transform 1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_125
timestamp 1698175906
transform 1 0 15344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_131
timestamp 1698175906
transform 1 0 16016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_135
timestamp 1698175906
transform 1 0 16464 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_151
timestamp 1698175906
transform 1 0 18256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_159
timestamp 1698175906
transform 1 0 19152 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_163
timestamp 1698175906
transform 1 0 19600 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_170
timestamp 1698175906
transform 1 0 20384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_96
timestamp 1698175906
transform 1 0 12096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_100
timestamp 1698175906
transform 1 0 12544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_102
timestamp 1698175906
transform 1 0 12768 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_150
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_152
timestamp 1698175906
transform 1 0 18368 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_183
timestamp 1698175906
transform 1 0 21840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_193
timestamp 1698175906
transform 1 0 22960 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_202
timestamp 1698175906
transform 1 0 23968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_218
timestamp 1698175906
transform 1 0 25760 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_250
timestamp 1698175906
transform 1 0 29344 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_266
timestamp 1698175906
transform 1 0 31136 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698175906
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698175906
transform 1 0 14000 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_143
timestamp 1698175906
transform 1 0 17360 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_182
timestamp 1698175906
transform 1 0 21728 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_215
timestamp 1698175906
transform 1 0 25424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_219
timestamp 1698175906
transform 1 0 25872 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_235
timestamp 1698175906
transform 1 0 27664 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_80
timestamp 1698175906
transform 1 0 10304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_84
timestamp 1698175906
transform 1 0 10752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_86
timestamp 1698175906
transform 1 0 10976 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_116
timestamp 1698175906
transform 1 0 14336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_118
timestamp 1698175906
transform 1 0 14560 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_146
timestamp 1698175906
transform 1 0 17696 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_154
timestamp 1698175906
transform 1 0 18592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_184
timestamp 1698175906
transform 1 0 21952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_188
timestamp 1698175906
transform 1 0 22400 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_115
timestamp 1698175906
transform 1 0 14224 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_118
timestamp 1698175906
transform 1 0 14560 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_150
timestamp 1698175906
transform 1 0 18144 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_166
timestamp 1698175906
transform 1 0 19936 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698175906
transform 1 0 19824 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_203
timestamp 1698175906
transform 1 0 24080 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_237
timestamp 1698175906
transform 1 0 27888 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 18592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_108
timestamp 1698175906
transform 1 0 13440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 4480 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 4480 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform -1 0 21616 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 4480 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 4480 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 16912 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 16576 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 24976 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 20384 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 4480 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform 1 0 21616 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 23520 41200 23632 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 41200 16800 42000 16912 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 21504 41200 21616 42000 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 19656 22736 19656 22736 0 _000_
rlabel metal2 24248 18872 24248 18872 0 _001_
rlabel metal2 22624 26936 22624 26936 0 _002_
rlabel metal2 24024 23520 24024 23520 0 _003_
rlabel metal2 24136 21952 24136 21952 0 _004_
rlabel metal3 13440 21784 13440 21784 0 _005_
rlabel metal2 26152 19264 26152 19264 0 _006_
rlabel metal2 12824 16128 12824 16128 0 _007_
rlabel metal2 12152 17976 12152 17976 0 _008_
rlabel metal3 14112 25704 14112 25704 0 _009_
rlabel metal2 18088 13048 18088 13048 0 _010_
rlabel metal2 15064 27384 15064 27384 0 _011_
rlabel metal2 13832 27216 13832 27216 0 _012_
rlabel metal2 15848 22568 15848 22568 0 _013_
rlabel metal2 13944 22456 13944 22456 0 _014_
rlabel metal2 26488 18032 26488 18032 0 _015_
rlabel metal2 20776 26656 20776 26656 0 _016_
rlabel metal2 18424 26908 18424 26908 0 _017_
rlabel metal2 19208 15484 19208 15484 0 _018_
rlabel metal2 22120 22064 22120 22064 0 _019_
rlabel metal2 24472 16744 24472 16744 0 _020_
rlabel metal2 11816 18760 11816 18760 0 _021_
rlabel metal2 14728 15792 14728 15792 0 _022_
rlabel metal2 26488 16520 26488 16520 0 _023_
rlabel metal2 14728 19656 14728 19656 0 _024_
rlabel metal2 19880 22792 19880 22792 0 _025_
rlabel metal2 17640 19712 17640 19712 0 _026_
rlabel metal2 27160 18816 27160 18816 0 _027_
rlabel metal2 16576 27608 16576 27608 0 _028_
rlabel metal2 14952 24640 14952 24640 0 _029_
rlabel metal3 23184 26264 23184 26264 0 _030_
rlabel metal3 25144 23016 25144 23016 0 _031_
rlabel metal2 24472 22288 24472 22288 0 _032_
rlabel metal2 14840 21896 14840 21896 0 _033_
rlabel metal2 15064 21952 15064 21952 0 _034_
rlabel metal2 15792 19432 15792 19432 0 _035_
rlabel metal2 28952 19432 28952 19432 0 _036_
rlabel metal2 26040 18816 26040 18816 0 _037_
rlabel metal2 14056 18816 14056 18816 0 _038_
rlabel metal2 14280 16576 14280 16576 0 _039_
rlabel metal3 14504 25368 14504 25368 0 _040_
rlabel metal2 15400 18704 15400 18704 0 _041_
rlabel metal2 14616 18592 14616 18592 0 _042_
rlabel metal2 14616 25368 14616 25368 0 _043_
rlabel metal2 17864 13944 17864 13944 0 _044_
rlabel metal2 17976 16268 17976 16268 0 _045_
rlabel metal2 16072 26488 16072 26488 0 _046_
rlabel metal2 15456 27832 15456 27832 0 _047_
rlabel metal2 16408 22120 16408 22120 0 _048_
rlabel metal2 17416 22400 17416 22400 0 _049_
rlabel metal2 14168 22960 14168 22960 0 _050_
rlabel metal2 14280 23016 14280 23016 0 _051_
rlabel metal2 27720 17360 27720 17360 0 _052_
rlabel metal2 25032 18200 25032 18200 0 _053_
rlabel metal2 20832 18536 20832 18536 0 _054_
rlabel metal3 24416 18424 24416 18424 0 _055_
rlabel metal3 19376 19208 19376 19208 0 _056_
rlabel metal2 17976 19936 17976 19936 0 _057_
rlabel metal2 21448 17696 21448 17696 0 _058_
rlabel metal2 21728 17528 21728 17528 0 _059_
rlabel metal2 21616 17752 21616 17752 0 _060_
rlabel metal3 20048 23800 20048 23800 0 _061_
rlabel metal2 19208 17584 19208 17584 0 _062_
rlabel metal3 17248 26264 17248 26264 0 _063_
rlabel metal2 21112 26600 21112 26600 0 _064_
rlabel metal2 17808 20104 17808 20104 0 _065_
rlabel metal2 20776 24976 20776 24976 0 _066_
rlabel metal3 15568 27832 15568 27832 0 _067_
rlabel metal3 22176 14280 22176 14280 0 _068_
rlabel metal2 21448 17024 21448 17024 0 _069_
rlabel metal2 18536 26376 18536 26376 0 _070_
rlabel metal3 24528 17528 24528 17528 0 _071_
rlabel metal2 19208 26208 19208 26208 0 _072_
rlabel metal3 17752 17640 17752 17640 0 _073_
rlabel metal2 23912 21896 23912 21896 0 _074_
rlabel metal2 19544 18536 19544 18536 0 _075_
rlabel metal2 18424 17304 18424 17304 0 _076_
rlabel metal3 18984 15400 18984 15400 0 _077_
rlabel metal2 19824 15288 19824 15288 0 _078_
rlabel metal2 22456 15680 22456 15680 0 _079_
rlabel metal2 20104 15344 20104 15344 0 _080_
rlabel metal2 18648 20720 18648 20720 0 _081_
rlabel metal2 15064 20272 15064 20272 0 _082_
rlabel metal2 24248 15736 24248 15736 0 _083_
rlabel metal3 16856 17640 16856 17640 0 _084_
rlabel metal2 17360 16744 17360 16744 0 _085_
rlabel metal3 15960 19320 15960 19320 0 _086_
rlabel metal3 20608 17752 20608 17752 0 _087_
rlabel metal2 15512 24752 15512 24752 0 _088_
rlabel metal2 15960 19544 15960 19544 0 _089_
rlabel metal2 14728 17136 14728 17136 0 _090_
rlabel metal2 15624 16520 15624 16520 0 _091_
rlabel metal3 23520 16968 23520 16968 0 _092_
rlabel metal3 22064 19208 22064 19208 0 _093_
rlabel metal2 27384 18312 27384 18312 0 _094_
rlabel metal2 26936 16856 26936 16856 0 _095_
rlabel metal2 19880 21616 19880 21616 0 _096_
rlabel metal2 17976 17976 17976 17976 0 _097_
rlabel metal2 19656 21952 19656 21952 0 _098_
rlabel metal3 2478 26936 2478 26936 0 clk
rlabel metal2 22680 20440 22680 20440 0 clknet_0_clk
rlabel metal2 13608 22736 13608 22736 0 clknet_1_0__leaf_clk
rlabel metal2 22232 27440 22232 27440 0 clknet_1_1__leaf_clk
rlabel metal2 21784 14504 21784 14504 0 dut18.count\[0\]
rlabel metal2 22400 16072 22400 16072 0 dut18.count\[1\]
rlabel metal2 13944 19152 13944 19152 0 dut18.count\[2\]
rlabel metal2 18760 15624 18760 15624 0 dut18.count\[3\]
rlabel metal2 21224 38024 21224 38024 0 net1
rlabel metal2 4312 16296 4312 16296 0 net10
rlabel metal3 6356 22344 6356 22344 0 net11
rlabel metal2 13720 23072 13720 23072 0 net12
rlabel metal2 28616 19936 28616 19936 0 net13
rlabel metal3 6356 23912 6356 23912 0 net14
rlabel metal2 37912 23184 37912 23184 0 net15
rlabel metal3 16744 27160 16744 27160 0 net16
rlabel metal2 15904 31920 15904 31920 0 net17
rlabel metal3 31920 23184 31920 23184 0 net18
rlabel metal2 24696 26656 24696 26656 0 net19
rlabel metal3 6356 19208 6356 19208 0 net2
rlabel metal2 27384 19152 27384 19152 0 net20
rlabel metal2 28616 16520 28616 16520 0 net21
rlabel metal2 20216 15204 20216 15204 0 net22
rlabel metal2 19656 38024 19656 38024 0 net23
rlabel metal2 4312 15344 4312 15344 0 net24
rlabel metal2 21448 27328 21448 27328 0 net25
rlabel metal2 21672 24472 21672 24472 0 net26
rlabel metal2 28616 17696 28616 17696 0 net3
rlabel metal2 17528 8568 17528 8568 0 net4
rlabel metal2 11256 27384 11256 27384 0 net5
rlabel metal2 25592 31864 25592 31864 0 net6
rlabel metal2 4088 15176 4088 15176 0 net7
rlabel metal2 21448 22932 21448 22932 0 net8
rlabel metal2 25032 32592 25032 32592 0 net9
rlabel metal2 22232 39746 22232 39746 0 segm[0]
rlabel metal3 1358 18872 1358 18872 0 segm[10]
rlabel metal2 40040 17640 40040 17640 0 segm[11]
rlabel metal2 18200 2058 18200 2058 0 segm[12]
rlabel metal3 1358 26264 1358 26264 0 segm[13]
rlabel metal2 24248 39354 24248 39354 0 segm[1]
rlabel metal3 1414 15512 1414 15512 0 segm[2]
rlabel metal2 20216 39186 20216 39186 0 segm[3]
rlabel metal2 23576 39746 23576 39746 0 segm[4]
rlabel metal3 1358 16184 1358 16184 0 segm[5]
rlabel metal3 1358 22232 1358 22232 0 segm[6]
rlabel metal3 1358 22904 1358 22904 0 segm[7]
rlabel metal2 40040 21112 40040 21112 0 segm[8]
rlabel metal3 1358 23576 1358 23576 0 segm[9]
rlabel metal2 40040 23800 40040 23800 0 sel[0]
rlabel metal2 16856 38962 16856 38962 0 sel[10]
rlabel metal2 16184 39746 16184 39746 0 sel[11]
rlabel metal3 40642 22904 40642 22904 0 sel[1]
rlabel metal2 24920 38962 24920 38962 0 sel[2]
rlabel metal2 40040 19656 40040 19656 0 sel[3]
rlabel metal2 40040 16800 40040 16800 0 sel[4]
rlabel metal3 21504 3640 21504 3640 0 sel[5]
rlabel metal2 19544 39746 19544 39746 0 sel[6]
rlabel metal3 1358 14840 1358 14840 0 sel[7]
rlabel metal2 20888 38962 20888 38962 0 sel[8]
rlabel metal2 21560 39354 21560 39354 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
