magic
tech gf180mcuD
magscale 1 5
timestamp 1699645711
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 9744 20600 9800 21000
rect 10416 20600 10472 21000
rect 12432 20600 12488 21000
rect 14448 20600 14504 21000
rect 7728 0 7784 400
rect 8400 0 8456 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12096 0 12152 400
rect 12432 0 12488 400
<< obsm2 >>
rect 966 20570 9714 20600
rect 9830 20570 10386 20600
rect 10502 20570 12402 20600
rect 12518 20570 14418 20600
rect 14534 20570 20146 20600
rect 966 430 20146 20570
rect 966 400 7698 430
rect 7814 400 8370 430
rect 8486 400 10050 430
rect 10166 400 10386 430
rect 10502 400 11394 430
rect 11510 400 11730 430
rect 11846 400 12066 430
rect 12182 400 12402 430
rect 12518 400 20146 430
<< metal3 >>
rect 0 13776 400 13832
rect 20600 13440 21000 13496
rect 0 13104 400 13160
rect 20600 13104 21000 13160
rect 20600 11760 21000 11816
rect 20600 11424 21000 11480
rect 20600 10416 21000 10472
rect 0 10080 400 10136
rect 0 9744 400 9800
rect 20600 9744 21000 9800
rect 0 9408 400 9464
rect 0 9072 400 9128
rect 20600 9072 21000 9128
rect 0 8400 400 8456
rect 20600 5712 21000 5768
<< obsm3 >>
rect 400 13862 20600 19222
rect 430 13746 20600 13862
rect 400 13526 20600 13746
rect 400 13410 20570 13526
rect 400 13190 20600 13410
rect 430 13074 20570 13190
rect 400 11846 20600 13074
rect 400 11730 20570 11846
rect 400 11510 20600 11730
rect 400 11394 20570 11510
rect 400 10502 20600 11394
rect 400 10386 20570 10502
rect 400 10166 20600 10386
rect 430 10050 20600 10166
rect 400 9830 20600 10050
rect 430 9714 20570 9830
rect 400 9494 20600 9714
rect 430 9378 20600 9494
rect 400 9158 20600 9378
rect 430 9042 20570 9158
rect 400 8486 20600 9042
rect 430 8370 20600 8486
rect 400 5798 20600 8370
rect 400 5682 20570 5798
rect 400 1554 20600 5682
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 11942 10145 12026 11359
<< labels >>
rlabel metal3 s 0 13776 400 13832 6 clk
port 1 nsew signal input
rlabel metal2 s 14448 20600 14504 21000 6 segm[0]
port 2 nsew signal output
rlabel metal3 s 0 13104 400 13160 6 segm[10]
port 3 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 segm[11]
port 4 nsew signal output
rlabel metal3 s 20600 11424 21000 11480 6 segm[12]
port 5 nsew signal output
rlabel metal2 s 12432 20600 12488 21000 6 segm[13]
port 6 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 segm[2]
port 8 nsew signal output
rlabel metal3 s 20600 5712 21000 5768 6 segm[3]
port 9 nsew signal output
rlabel metal2 s 11424 0 11480 400 6 segm[4]
port 10 nsew signal output
rlabel metal3 s 0 10080 400 10136 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 20600 9744 21000 9800 6 segm[6]
port 12 nsew signal output
rlabel metal2 s 10416 20600 10472 21000 6 segm[7]
port 13 nsew signal output
rlabel metal3 s 20600 13440 21000 13496 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 20600 13104 21000 13160 6 segm[9]
port 15 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 sel[0]
port 16 nsew signal output
rlabel metal2 s 9744 20600 9800 21000 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 sel[11]
port 18 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 sel[1]
port 19 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 sel[2]
port 20 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 sel[3]
port 21 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 sel[4]
port 22 nsew signal output
rlabel metal2 s 7728 0 7784 400 6 sel[5]
port 23 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 sel[6]
port 24 nsew signal output
rlabel metal2 s 10080 0 10136 400 6 sel[7]
port 25 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 sel[8]
port 26 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 483526
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita40/runs/23_11_10_13_46/results/signoff/ita40.magic.gds
string GDS_START 155706
<< end >>

