magic
tech gf180mcuD
magscale 1 5
timestamp 1699641242
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 8400 20600 8456 21000
rect 9072 20600 9128 21000
rect 9408 20600 9464 21000
rect 10416 20600 10472 21000
rect 11088 20600 11144 21000
rect 11760 20600 11816 21000
rect 12096 20600 12152 21000
rect 3696 0 3752 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 12768 0 12824 400
<< obsm2 >>
rect 966 20570 8370 20600
rect 8486 20570 9042 20600
rect 9158 20570 9378 20600
rect 9494 20570 10386 20600
rect 10502 20570 11058 20600
rect 11174 20570 11730 20600
rect 11846 20570 12066 20600
rect 12182 20570 20146 20600
rect 966 430 20146 20570
rect 966 400 3666 430
rect 3782 400 10722 430
rect 10838 400 11058 430
rect 11174 400 12738 430
rect 12854 400 20146 430
<< metal3 >>
rect 20600 18480 21000 18536
rect 0 13776 400 13832
rect 20600 13440 21000 13496
rect 20600 13104 21000 13160
rect 20600 12768 21000 12824
rect 0 12432 400 12488
rect 20600 12432 21000 12488
rect 20600 10752 21000 10808
rect 0 10416 400 10472
rect 20600 10416 21000 10472
rect 20600 10080 21000 10136
rect 0 9072 400 9128
rect 0 8736 400 8792
rect 20600 8736 21000 8792
rect 0 8400 400 8456
rect 20600 8400 21000 8456
<< obsm3 >>
rect 400 18566 20600 19222
rect 400 18450 20570 18566
rect 400 13862 20600 18450
rect 430 13746 20600 13862
rect 400 13526 20600 13746
rect 400 13410 20570 13526
rect 400 13190 20600 13410
rect 400 13074 20570 13190
rect 400 12854 20600 13074
rect 400 12738 20570 12854
rect 400 12518 20600 12738
rect 430 12402 20570 12518
rect 400 10838 20600 12402
rect 400 10722 20570 10838
rect 400 10502 20600 10722
rect 430 10386 20570 10502
rect 400 10166 20600 10386
rect 400 10050 20570 10166
rect 400 9158 20600 10050
rect 430 9042 20600 9158
rect 400 8822 20600 9042
rect 430 8706 20570 8822
rect 400 8486 20600 8706
rect 430 8370 20570 8486
rect 400 1554 20600 8370
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 8022 8745 8050 9623
<< labels >>
rlabel metal3 s 0 13776 400 13832 6 clk
port 1 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 segm[0]
port 2 nsew signal output
rlabel metal2 s 11088 20600 11144 21000 6 segm[10]
port 3 nsew signal output
rlabel metal3 s 20600 10752 21000 10808 6 segm[11]
port 4 nsew signal output
rlabel metal2 s 8400 20600 8456 21000 6 segm[12]
port 5 nsew signal output
rlabel metal2 s 10752 0 10808 400 6 segm[13]
port 6 nsew signal output
rlabel metal3 s 20600 13440 21000 13496 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 segm[2]
port 8 nsew signal output
rlabel metal2 s 9408 20600 9464 21000 6 segm[3]
port 9 nsew signal output
rlabel metal3 s 20600 12768 21000 12824 6 segm[4]
port 10 nsew signal output
rlabel metal3 s 20600 18480 21000 18536 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 segm[6]
port 12 nsew signal output
rlabel metal3 s 20600 10080 21000 10136 6 segm[7]
port 13 nsew signal output
rlabel metal2 s 12096 20600 12152 21000 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 segm[9]
port 15 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 sel[0]
port 16 nsew signal output
rlabel metal2 s 11088 0 11144 400 6 sel[10]
port 17 nsew signal output
rlabel metal2 s 12768 0 12824 400 6 sel[11]
port 18 nsew signal output
rlabel metal2 s 10416 20600 10472 21000 6 sel[1]
port 19 nsew signal output
rlabel metal3 s 20600 8736 21000 8792 6 sel[2]
port 20 nsew signal output
rlabel metal2 s 11760 20600 11816 21000 6 sel[3]
port 21 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 sel[4]
port 22 nsew signal output
rlabel metal3 s 20600 13104 21000 13160 6 sel[5]
port 23 nsew signal output
rlabel metal2 s 9072 20600 9128 21000 6 sel[6]
port 24 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 sel[7]
port 25 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 sel[8]
port 26 nsew signal output
rlabel metal3 s 20600 8400 21000 8456 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 489676
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita2/runs/23_11_10_12_32/results/signoff/ita2.magic.gds
string GDS_START 172476
<< end >>

