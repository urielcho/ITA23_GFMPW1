magic
tech gf180mcuD
magscale 1 10
timestamp 1699642593
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 22094 38274 22146 38286
rect 22094 38210 22146 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 17938 37998 17950 38050
rect 18002 37998 18014 38050
rect 21186 37998 21198 38050
rect 21250 37998 21262 38050
rect 24994 37998 25006 38050
rect 25058 37998 25070 38050
rect 27470 37938 27522 37950
rect 27470 37874 27522 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18510 37490 18562 37502
rect 18510 37426 18562 37438
rect 21422 37490 21474 37502
rect 21422 37426 21474 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 17602 37214 17614 37266
rect 17666 37214 17678 37266
rect 20626 37214 20638 37266
rect 20690 37214 20702 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 18062 36706 18114 36718
rect 18062 36642 18114 36654
rect 17378 36430 17390 36482
rect 17442 36430 17454 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 17378 28702 17390 28754
rect 17442 28702 17454 28754
rect 18510 28642 18562 28654
rect 14578 28590 14590 28642
rect 14642 28590 14654 28642
rect 18510 28578 18562 28590
rect 21758 28642 21810 28654
rect 21758 28578 21810 28590
rect 17726 28530 17778 28542
rect 15250 28478 15262 28530
rect 15314 28478 15326 28530
rect 18050 28478 18062 28530
rect 18114 28478 18126 28530
rect 17726 28466 17778 28478
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 15934 28082 15986 28094
rect 15934 28018 15986 28030
rect 16718 28082 16770 28094
rect 16718 28018 16770 28030
rect 17390 28082 17442 28094
rect 17714 28030 17726 28082
rect 17778 28030 17790 28082
rect 17390 28018 17442 28030
rect 16158 27970 16210 27982
rect 16158 27906 16210 27918
rect 16270 27858 16322 27870
rect 16270 27794 16322 27806
rect 16494 27858 16546 27870
rect 16494 27794 16546 27806
rect 16830 27858 16882 27870
rect 18610 27806 18622 27858
rect 18674 27806 18686 27858
rect 21746 27806 21758 27858
rect 21810 27806 21822 27858
rect 16830 27794 16882 27806
rect 25342 27746 25394 27758
rect 19282 27694 19294 27746
rect 19346 27694 19358 27746
rect 21410 27694 21422 27746
rect 21474 27694 21486 27746
rect 22530 27694 22542 27746
rect 22594 27694 22606 27746
rect 24658 27694 24670 27746
rect 24722 27694 24734 27746
rect 25342 27682 25394 27694
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 25454 27298 25506 27310
rect 25454 27234 25506 27246
rect 40014 27186 40066 27198
rect 20626 27134 20638 27186
rect 20690 27134 20702 27186
rect 25106 27134 25118 27186
rect 25170 27134 25182 27186
rect 40014 27122 40066 27134
rect 17826 27022 17838 27074
rect 17890 27022 17902 27074
rect 22306 27022 22318 27074
rect 22370 27022 22382 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 21422 26962 21474 26974
rect 18498 26910 18510 26962
rect 18562 26910 18574 26962
rect 21422 26898 21474 26910
rect 21534 26962 21586 26974
rect 25566 26962 25618 26974
rect 22978 26910 22990 26962
rect 23042 26910 23054 26962
rect 21534 26898 21586 26910
rect 25566 26898 25618 26910
rect 21198 26850 21250 26862
rect 21198 26786 21250 26798
rect 26014 26850 26066 26862
rect 26014 26786 26066 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 19070 26514 19122 26526
rect 17378 26462 17390 26514
rect 17442 26462 17454 26514
rect 19070 26450 19122 26462
rect 19742 26514 19794 26526
rect 19742 26450 19794 26462
rect 20526 26514 20578 26526
rect 20526 26450 20578 26462
rect 21422 26514 21474 26526
rect 21422 26450 21474 26462
rect 22654 26514 22706 26526
rect 22654 26450 22706 26462
rect 23326 26514 23378 26526
rect 23326 26450 23378 26462
rect 23438 26514 23490 26526
rect 23438 26450 23490 26462
rect 23550 26514 23602 26526
rect 23550 26450 23602 26462
rect 24334 26514 24386 26526
rect 24334 26450 24386 26462
rect 24446 26514 24498 26526
rect 24446 26450 24498 26462
rect 24558 26514 24610 26526
rect 24558 26450 24610 26462
rect 18958 26402 19010 26414
rect 18958 26338 19010 26350
rect 17726 26290 17778 26302
rect 4274 26238 4286 26290
rect 4338 26238 4350 26290
rect 15586 26238 15598 26290
rect 15650 26238 15662 26290
rect 17726 26226 17778 26238
rect 19518 26290 19570 26302
rect 19518 26226 19570 26238
rect 20190 26290 20242 26302
rect 20190 26226 20242 26238
rect 20414 26290 20466 26302
rect 20414 26226 20466 26238
rect 20638 26290 20690 26302
rect 20638 26226 20690 26238
rect 21086 26290 21138 26302
rect 21086 26226 21138 26238
rect 22542 26290 22594 26302
rect 22542 26226 22594 26238
rect 23102 26290 23154 26302
rect 23102 26226 23154 26238
rect 23214 26290 23266 26302
rect 23214 26226 23266 26238
rect 24110 26290 24162 26302
rect 24110 26226 24162 26238
rect 24222 26290 24274 26302
rect 25442 26238 25454 26290
rect 25506 26238 25518 26290
rect 24222 26226 24274 26238
rect 16046 26178 16098 26190
rect 12674 26126 12686 26178
rect 12738 26126 12750 26178
rect 14802 26126 14814 26178
rect 14866 26126 14878 26178
rect 16046 26114 16098 26126
rect 16830 26178 16882 26190
rect 16830 26114 16882 26126
rect 19630 26178 19682 26190
rect 26226 26126 26238 26178
rect 26290 26126 26302 26178
rect 28354 26126 28366 26178
rect 28418 26126 28430 26178
rect 19630 26114 19682 26126
rect 1934 26066 1986 26078
rect 1934 26002 1986 26014
rect 19182 26066 19234 26078
rect 19182 26002 19234 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 16830 25618 16882 25630
rect 2034 25566 2046 25618
rect 2098 25566 2110 25618
rect 16370 25566 16382 25618
rect 16434 25566 16446 25618
rect 16830 25554 16882 25566
rect 17502 25618 17554 25630
rect 17502 25554 17554 25566
rect 26014 25618 26066 25630
rect 26014 25554 26066 25566
rect 26574 25506 26626 25518
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 13570 25454 13582 25506
rect 13634 25454 13646 25506
rect 17042 25454 17054 25506
rect 17106 25454 17118 25506
rect 26574 25442 26626 25454
rect 27022 25506 27074 25518
rect 27022 25442 27074 25454
rect 27358 25506 27410 25518
rect 27358 25442 27410 25454
rect 27806 25506 27858 25518
rect 27806 25442 27858 25454
rect 16718 25394 16770 25406
rect 14242 25342 14254 25394
rect 14306 25342 14318 25394
rect 16718 25330 16770 25342
rect 27246 25394 27298 25406
rect 27246 25330 27298 25342
rect 25118 25282 25170 25294
rect 25118 25218 25170 25230
rect 25902 25282 25954 25294
rect 25902 25218 25954 25230
rect 26126 25282 26178 25294
rect 26126 25218 26178 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 14590 24946 14642 24958
rect 14590 24882 14642 24894
rect 16158 24946 16210 24958
rect 16158 24882 16210 24894
rect 17614 24946 17666 24958
rect 17614 24882 17666 24894
rect 18398 24946 18450 24958
rect 18398 24882 18450 24894
rect 22542 24946 22594 24958
rect 22542 24882 22594 24894
rect 16270 24834 16322 24846
rect 16270 24770 16322 24782
rect 18286 24834 18338 24846
rect 18286 24770 18338 24782
rect 21310 24834 21362 24846
rect 21310 24770 21362 24782
rect 22318 24834 22370 24846
rect 22318 24770 22370 24782
rect 17390 24722 17442 24734
rect 15922 24670 15934 24722
rect 15986 24670 15998 24722
rect 17390 24658 17442 24670
rect 18062 24722 18114 24734
rect 18062 24658 18114 24670
rect 18622 24722 18674 24734
rect 21198 24722 21250 24734
rect 20738 24670 20750 24722
rect 20802 24670 20814 24722
rect 18622 24658 18674 24670
rect 21198 24658 21250 24670
rect 22206 24722 22258 24734
rect 37650 24670 37662 24722
rect 37714 24670 37726 24722
rect 22206 24658 22258 24670
rect 14702 24610 14754 24622
rect 14702 24546 14754 24558
rect 17502 24610 17554 24622
rect 17502 24546 17554 24558
rect 20974 24498 21026 24510
rect 20974 24434 21026 24446
rect 40014 24498 40066 24510
rect 40014 24434 40066 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 16270 24162 16322 24174
rect 16270 24098 16322 24110
rect 16606 24162 16658 24174
rect 16606 24098 16658 24110
rect 18958 24162 19010 24174
rect 18958 24098 19010 24110
rect 28578 23998 28590 24050
rect 28642 23998 28654 24050
rect 17602 23886 17614 23938
rect 17666 23886 17678 23938
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 16830 23826 16882 23838
rect 18622 23826 18674 23838
rect 17826 23774 17838 23826
rect 17890 23774 17902 23826
rect 16830 23762 16882 23774
rect 18622 23762 18674 23774
rect 18846 23826 18898 23838
rect 18846 23762 18898 23774
rect 22542 23826 22594 23838
rect 23202 23774 23214 23826
rect 23266 23774 23278 23826
rect 26450 23774 26462 23826
rect 26514 23774 26526 23826
rect 22542 23762 22594 23774
rect 22206 23714 22258 23726
rect 22206 23650 22258 23662
rect 22430 23714 22482 23726
rect 22430 23650 22482 23662
rect 22878 23714 22930 23726
rect 22878 23650 22930 23662
rect 25342 23714 25394 23726
rect 25342 23650 25394 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 16382 23378 16434 23390
rect 16382 23314 16434 23326
rect 17726 23378 17778 23390
rect 18846 23378 18898 23390
rect 18050 23326 18062 23378
rect 18114 23326 18126 23378
rect 17726 23314 17778 23326
rect 18846 23314 18898 23326
rect 19182 23378 19234 23390
rect 19182 23314 19234 23326
rect 23774 23378 23826 23390
rect 23774 23314 23826 23326
rect 26350 23378 26402 23390
rect 26350 23314 26402 23326
rect 27358 23378 27410 23390
rect 27358 23314 27410 23326
rect 27918 23378 27970 23390
rect 27918 23314 27970 23326
rect 18622 23266 18674 23278
rect 18622 23202 18674 23214
rect 19070 23266 19122 23278
rect 19070 23202 19122 23214
rect 19630 23266 19682 23278
rect 19630 23202 19682 23214
rect 23550 23266 23602 23278
rect 23550 23202 23602 23214
rect 23998 23266 24050 23278
rect 23998 23202 24050 23214
rect 27470 23266 27522 23278
rect 27470 23202 27522 23214
rect 16046 23154 16098 23166
rect 16046 23090 16098 23102
rect 19518 23154 19570 23166
rect 19518 23090 19570 23102
rect 19854 23154 19906 23166
rect 19854 23090 19906 23102
rect 20078 23154 20130 23166
rect 26238 23154 26290 23166
rect 20402 23102 20414 23154
rect 20466 23102 20478 23154
rect 21074 23102 21086 23154
rect 21138 23102 21150 23154
rect 20078 23090 20130 23102
rect 26238 23090 26290 23102
rect 26462 23154 26514 23166
rect 26462 23090 26514 23102
rect 26910 23154 26962 23166
rect 26910 23090 26962 23102
rect 27134 23154 27186 23166
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 27134 23090 27186 23102
rect 15374 23042 15426 23054
rect 24446 23042 24498 23054
rect 23202 22990 23214 23042
rect 23266 22990 23278 23042
rect 15374 22978 15426 22990
rect 24446 22978 24498 22990
rect 15486 22930 15538 22942
rect 15486 22866 15538 22878
rect 23662 22930 23714 22942
rect 23662 22866 23714 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 13582 22482 13634 22494
rect 12898 22430 12910 22482
rect 12962 22430 12974 22482
rect 13582 22418 13634 22430
rect 14030 22482 14082 22494
rect 14030 22418 14082 22430
rect 27022 22482 27074 22494
rect 27022 22418 27074 22430
rect 40014 22482 40066 22494
rect 40014 22418 40066 22430
rect 15486 22370 15538 22382
rect 10098 22318 10110 22370
rect 10162 22318 10174 22370
rect 14578 22318 14590 22370
rect 14642 22318 14654 22370
rect 15486 22306 15538 22318
rect 15934 22370 15986 22382
rect 15934 22306 15986 22318
rect 16494 22370 16546 22382
rect 16494 22306 16546 22318
rect 16830 22370 16882 22382
rect 16830 22306 16882 22318
rect 17054 22370 17106 22382
rect 17054 22306 17106 22318
rect 17726 22370 17778 22382
rect 26798 22370 26850 22382
rect 21970 22318 21982 22370
rect 22034 22318 22046 22370
rect 37874 22318 37886 22370
rect 37938 22318 37950 22370
rect 17726 22306 17778 22318
rect 26798 22306 26850 22318
rect 10770 22206 10782 22258
rect 10834 22206 10846 22258
rect 25778 22206 25790 22258
rect 25842 22206 25854 22258
rect 14142 22146 14194 22158
rect 15598 22146 15650 22158
rect 14802 22094 14814 22146
rect 14866 22094 14878 22146
rect 14142 22082 14194 22094
rect 15598 22082 15650 22094
rect 16718 22146 16770 22158
rect 16718 22082 16770 22094
rect 17390 22146 17442 22158
rect 17390 22082 17442 22094
rect 17614 22146 17666 22158
rect 17614 22082 17666 22094
rect 18846 22146 18898 22158
rect 27134 22146 27186 22158
rect 19170 22094 19182 22146
rect 19234 22094 19246 22146
rect 18846 22082 18898 22094
rect 27134 22082 27186 22094
rect 27358 22146 27410 22158
rect 27358 22082 27410 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14254 21810 14306 21822
rect 14254 21746 14306 21758
rect 15038 21810 15090 21822
rect 15038 21746 15090 21758
rect 17614 21810 17666 21822
rect 17614 21746 17666 21758
rect 24110 21810 24162 21822
rect 24110 21746 24162 21758
rect 15822 21698 15874 21710
rect 11666 21646 11678 21698
rect 11730 21646 11742 21698
rect 15362 21646 15374 21698
rect 15426 21646 15438 21698
rect 15822 21634 15874 21646
rect 24334 21698 24386 21710
rect 24334 21634 24386 21646
rect 15710 21586 15762 21598
rect 10994 21534 11006 21586
rect 11058 21534 11070 21586
rect 15710 21522 15762 21534
rect 15934 21586 15986 21598
rect 16258 21534 16270 21586
rect 16322 21534 16334 21586
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 18162 21534 18174 21586
rect 18226 21534 18238 21586
rect 23874 21534 23886 21586
rect 23938 21534 23950 21586
rect 25778 21534 25790 21586
rect 25842 21534 25854 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 15934 21522 15986 21534
rect 23998 21474 24050 21486
rect 13794 21422 13806 21474
rect 13858 21422 13870 21474
rect 20290 21422 20302 21474
rect 20354 21422 20366 21474
rect 23998 21410 24050 21422
rect 25454 21474 25506 21486
rect 40014 21474 40066 21486
rect 26562 21422 26574 21474
rect 26626 21422 26638 21474
rect 28690 21422 28702 21474
rect 28754 21422 28766 21474
rect 25454 21410 25506 21422
rect 40014 21410 40066 21422
rect 17502 21362 17554 21374
rect 17502 21298 17554 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 26798 21026 26850 21038
rect 14690 20974 14702 21026
rect 14754 21023 14766 21026
rect 14914 21023 14926 21026
rect 14754 20977 14926 21023
rect 14754 20974 14766 20977
rect 14914 20974 14926 20977
rect 14978 20974 14990 21026
rect 26798 20962 26850 20974
rect 14926 20914 14978 20926
rect 14926 20850 14978 20862
rect 17950 20914 18002 20926
rect 27358 20914 27410 20926
rect 23650 20862 23662 20914
rect 23714 20862 23726 20914
rect 25778 20862 25790 20914
rect 25842 20862 25854 20914
rect 17950 20850 18002 20862
rect 27358 20850 27410 20862
rect 15486 20802 15538 20814
rect 16158 20802 16210 20814
rect 15810 20750 15822 20802
rect 15874 20750 15886 20802
rect 15486 20738 15538 20750
rect 16158 20738 16210 20750
rect 18846 20802 18898 20814
rect 19854 20802 19906 20814
rect 19618 20750 19630 20802
rect 19682 20750 19694 20802
rect 18846 20738 18898 20750
rect 19854 20738 19906 20750
rect 20190 20802 20242 20814
rect 20190 20738 20242 20750
rect 21534 20802 21586 20814
rect 21534 20738 21586 20750
rect 22206 20802 22258 20814
rect 22866 20750 22878 20802
rect 22930 20750 22942 20802
rect 22206 20738 22258 20750
rect 20078 20690 20130 20702
rect 26238 20690 26290 20702
rect 16706 20638 16718 20690
rect 16770 20638 16782 20690
rect 18498 20638 18510 20690
rect 18562 20638 18574 20690
rect 21858 20638 21870 20690
rect 21922 20638 21934 20690
rect 20078 20626 20130 20638
rect 26238 20626 26290 20638
rect 26350 20690 26402 20702
rect 26350 20626 26402 20638
rect 26686 20690 26738 20702
rect 26686 20626 26738 20638
rect 26798 20690 26850 20702
rect 26798 20626 26850 20638
rect 16046 20578 16098 20590
rect 16046 20514 16098 20526
rect 16382 20578 16434 20590
rect 16382 20514 16434 20526
rect 18174 20578 18226 20590
rect 19966 20578 20018 20590
rect 26014 20578 26066 20590
rect 19170 20526 19182 20578
rect 19234 20526 19246 20578
rect 22530 20526 22542 20578
rect 22594 20526 22606 20578
rect 18174 20514 18226 20526
rect 19966 20514 20018 20526
rect 26014 20514 26066 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 15150 20242 15202 20254
rect 15150 20178 15202 20190
rect 19070 20242 19122 20254
rect 19070 20178 19122 20190
rect 19966 20242 20018 20254
rect 19966 20178 20018 20190
rect 25902 20242 25954 20254
rect 25902 20178 25954 20190
rect 17726 20130 17778 20142
rect 15922 20078 15934 20130
rect 15986 20078 15998 20130
rect 17726 20066 17778 20078
rect 18510 20130 18562 20142
rect 18510 20066 18562 20078
rect 18622 20130 18674 20142
rect 18622 20066 18674 20078
rect 19406 20130 19458 20142
rect 19406 20066 19458 20078
rect 20526 20130 20578 20142
rect 20526 20066 20578 20078
rect 20638 20130 20690 20142
rect 20638 20066 20690 20078
rect 21534 20130 21586 20142
rect 21534 20066 21586 20078
rect 21758 20130 21810 20142
rect 21758 20066 21810 20078
rect 21982 20130 22034 20142
rect 21982 20066 22034 20078
rect 22094 20130 22146 20142
rect 22094 20066 22146 20078
rect 22318 20130 22370 20142
rect 22318 20066 22370 20078
rect 24334 20130 24386 20142
rect 25342 20130 25394 20142
rect 24658 20078 24670 20130
rect 24722 20078 24734 20130
rect 24334 20066 24386 20078
rect 25342 20066 25394 20078
rect 25790 20130 25842 20142
rect 25790 20066 25842 20078
rect 26126 20130 26178 20142
rect 26126 20066 26178 20078
rect 26350 20130 26402 20142
rect 26350 20066 26402 20078
rect 26574 20130 26626 20142
rect 26574 20066 26626 20078
rect 14814 20018 14866 20030
rect 17390 20018 17442 20030
rect 15586 19966 15598 20018
rect 15650 19966 15662 20018
rect 14814 19954 14866 19966
rect 17390 19954 17442 19966
rect 18286 20018 18338 20030
rect 18286 19954 18338 19966
rect 19294 20018 19346 20030
rect 19294 19954 19346 19966
rect 19518 20018 19570 20030
rect 19518 19954 19570 19966
rect 19742 20018 19794 20030
rect 19742 19954 19794 19966
rect 20078 20018 20130 20030
rect 20078 19954 20130 19966
rect 21422 20018 21474 20030
rect 25554 19966 25566 20018
rect 25618 19966 25630 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 21422 19954 21474 19966
rect 13806 19906 13858 19918
rect 15026 19854 15038 19906
rect 15090 19854 15102 19906
rect 16258 19854 16270 19906
rect 16322 19854 16334 19906
rect 13806 19842 13858 19854
rect 13918 19794 13970 19806
rect 13918 19730 13970 19742
rect 20526 19794 20578 19806
rect 20526 19730 20578 19742
rect 26238 19794 26290 19806
rect 26238 19730 26290 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 40014 19346 40066 19358
rect 15250 19294 15262 19346
rect 15314 19294 15326 19346
rect 24770 19294 24782 19346
rect 24834 19294 24846 19346
rect 28018 19294 28030 19346
rect 28082 19294 28094 19346
rect 40014 19282 40066 19294
rect 13470 19234 13522 19246
rect 13470 19170 13522 19182
rect 14478 19234 14530 19246
rect 14478 19170 14530 19182
rect 14702 19234 14754 19246
rect 21198 19234 21250 19246
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 14702 19170 14754 19182
rect 21198 19170 21250 19182
rect 21422 19234 21474 19246
rect 21422 19170 21474 19182
rect 21646 19234 21698 19246
rect 21646 19170 21698 19182
rect 21870 19234 21922 19246
rect 21870 19170 21922 19182
rect 22206 19234 22258 19246
rect 25218 19182 25230 19234
rect 25282 19182 25294 19234
rect 37650 19182 37662 19234
rect 37714 19182 37726 19234
rect 22206 19170 22258 19182
rect 24334 19122 24386 19134
rect 24546 19070 24558 19122
rect 24610 19070 24622 19122
rect 25890 19070 25902 19122
rect 25954 19070 25966 19122
rect 24334 19058 24386 19070
rect 14254 19010 14306 19022
rect 13794 18958 13806 19010
rect 13858 18958 13870 19010
rect 14254 18946 14306 18958
rect 14590 19010 14642 19022
rect 23662 19010 23714 19022
rect 22530 18958 22542 19010
rect 22594 18958 22606 19010
rect 14590 18946 14642 18958
rect 23662 18946 23714 18958
rect 23998 19010 24050 19022
rect 23998 18946 24050 18958
rect 24222 19010 24274 19022
rect 24222 18946 24274 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 14814 18674 14866 18686
rect 14814 18610 14866 18622
rect 19630 18674 19682 18686
rect 21310 18674 21362 18686
rect 19954 18622 19966 18674
rect 20018 18622 20030 18674
rect 19630 18610 19682 18622
rect 21310 18610 21362 18622
rect 15038 18562 15090 18574
rect 16830 18562 16882 18574
rect 15362 18510 15374 18562
rect 15426 18510 15438 18562
rect 15038 18498 15090 18510
rect 16830 18498 16882 18510
rect 17390 18562 17442 18574
rect 17390 18498 17442 18510
rect 17726 18562 17778 18574
rect 17726 18498 17778 18510
rect 18846 18562 18898 18574
rect 20974 18562 21026 18574
rect 20626 18510 20638 18562
rect 20690 18510 20702 18562
rect 18846 18498 18898 18510
rect 20974 18498 21026 18510
rect 21086 18562 21138 18574
rect 21086 18498 21138 18510
rect 14142 18450 14194 18462
rect 16046 18450 16098 18462
rect 4274 18398 4286 18450
rect 4338 18398 4350 18450
rect 10658 18398 10670 18450
rect 10722 18398 10734 18450
rect 15250 18398 15262 18450
rect 15314 18398 15326 18450
rect 14142 18386 14194 18398
rect 16046 18386 16098 18398
rect 16606 18450 16658 18462
rect 16606 18386 16658 18398
rect 18510 18450 18562 18462
rect 18510 18386 18562 18398
rect 20302 18450 20354 18462
rect 25330 18398 25342 18450
rect 25394 18398 25406 18450
rect 26002 18398 26014 18450
rect 26066 18398 26078 18450
rect 20302 18386 20354 18398
rect 13918 18338 13970 18350
rect 24670 18338 24722 18350
rect 11330 18286 11342 18338
rect 11394 18286 11406 18338
rect 13458 18286 13470 18338
rect 13522 18286 13534 18338
rect 15026 18286 15038 18338
rect 15090 18286 15102 18338
rect 16482 18286 16494 18338
rect 16546 18286 16558 18338
rect 18162 18286 18174 18338
rect 18226 18286 18238 18338
rect 28130 18286 28142 18338
rect 28194 18286 28206 18338
rect 13918 18274 13970 18286
rect 24670 18274 24722 18286
rect 1934 18226 1986 18238
rect 16270 18226 16322 18238
rect 14466 18174 14478 18226
rect 14530 18174 14542 18226
rect 1934 18162 1986 18174
rect 16270 18162 16322 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 14366 17890 14418 17902
rect 14366 17826 14418 17838
rect 14702 17890 14754 17902
rect 16494 17890 16546 17902
rect 15586 17838 15598 17890
rect 15650 17838 15662 17890
rect 14702 17826 14754 17838
rect 16494 17826 16546 17838
rect 19182 17890 19234 17902
rect 19182 17826 19234 17838
rect 13694 17778 13746 17790
rect 13694 17714 13746 17726
rect 18958 17778 19010 17790
rect 18958 17714 19010 17726
rect 15038 17666 15090 17678
rect 16718 17666 16770 17678
rect 15250 17614 15262 17666
rect 15314 17614 15326 17666
rect 15698 17614 15710 17666
rect 15762 17614 15774 17666
rect 16146 17614 16158 17666
rect 16210 17614 16222 17666
rect 15038 17602 15090 17614
rect 16718 17602 16770 17614
rect 18622 17666 18674 17678
rect 18622 17602 18674 17614
rect 19854 17666 19906 17678
rect 22306 17614 22318 17666
rect 22370 17614 22382 17666
rect 19854 17602 19906 17614
rect 14478 17554 14530 17566
rect 20190 17554 20242 17566
rect 17378 17502 17390 17554
rect 17442 17502 17454 17554
rect 14478 17490 14530 17502
rect 20190 17490 20242 17502
rect 22766 17554 22818 17566
rect 22766 17490 22818 17502
rect 15150 17442 15202 17454
rect 15150 17378 15202 17390
rect 17054 17442 17106 17454
rect 17054 17378 17106 17390
rect 18510 17442 18562 17454
rect 22878 17442 22930 17454
rect 19506 17390 19518 17442
rect 19570 17390 19582 17442
rect 18510 17378 18562 17390
rect 22878 17378 22930 17390
rect 22990 17442 23042 17454
rect 22990 17378 23042 17390
rect 23102 17442 23154 17454
rect 23102 17378 23154 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 21198 17106 21250 17118
rect 21198 17042 21250 17054
rect 21422 17106 21474 17118
rect 21422 17042 21474 17054
rect 22542 17106 22594 17118
rect 22542 17042 22594 17054
rect 23438 17106 23490 17118
rect 23438 17042 23490 17054
rect 23662 17106 23714 17118
rect 23662 17042 23714 17054
rect 21534 16994 21586 17006
rect 22654 16994 22706 17006
rect 13010 16942 13022 16994
rect 13074 16942 13086 16994
rect 21634 16942 21646 16994
rect 21698 16942 21710 16994
rect 21534 16930 21586 16942
rect 22654 16930 22706 16942
rect 23774 16994 23826 17006
rect 23774 16930 23826 16942
rect 14254 16882 14306 16894
rect 13682 16830 13694 16882
rect 13746 16830 13758 16882
rect 14254 16818 14306 16830
rect 22318 16882 22370 16894
rect 22978 16830 22990 16882
rect 23042 16830 23054 16882
rect 24210 16830 24222 16882
rect 24274 16830 24286 16882
rect 22318 16818 22370 16830
rect 22430 16770 22482 16782
rect 10882 16718 10894 16770
rect 10946 16718 10958 16770
rect 21970 16718 21982 16770
rect 22034 16718 22046 16770
rect 22430 16706 22482 16718
rect 23550 16770 23602 16782
rect 23550 16706 23602 16718
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 18062 16322 18114 16334
rect 18062 16258 18114 16270
rect 23986 16158 23998 16210
rect 24050 16158 24062 16210
rect 26114 16158 26126 16210
rect 26178 16158 26190 16210
rect 17278 16098 17330 16110
rect 17278 16034 17330 16046
rect 17502 16098 17554 16110
rect 17714 16046 17726 16098
rect 17778 16046 17790 16098
rect 19394 16046 19406 16098
rect 19458 16046 19470 16098
rect 23202 16046 23214 16098
rect 23266 16046 23278 16098
rect 17502 16034 17554 16046
rect 19170 15934 19182 15986
rect 19234 15934 19246 15986
rect 17614 15874 17666 15886
rect 17614 15810 17666 15822
rect 18174 15874 18226 15886
rect 18174 15810 18226 15822
rect 18286 15874 18338 15886
rect 18286 15810 18338 15822
rect 26574 15874 26626 15886
rect 26574 15810 26626 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 15038 15538 15090 15550
rect 15038 15474 15090 15486
rect 21086 15538 21138 15550
rect 21086 15474 21138 15486
rect 20078 15426 20130 15438
rect 12450 15374 12462 15426
rect 12514 15374 12526 15426
rect 17938 15374 17950 15426
rect 18002 15374 18014 15426
rect 22082 15374 22094 15426
rect 22146 15374 22158 15426
rect 20078 15362 20130 15374
rect 16382 15314 16434 15326
rect 11778 15262 11790 15314
rect 11842 15262 11854 15314
rect 16382 15250 16434 15262
rect 16606 15314 16658 15326
rect 18174 15314 18226 15326
rect 17602 15262 17614 15314
rect 17666 15262 17678 15314
rect 16606 15250 16658 15262
rect 18174 15250 18226 15262
rect 18510 15314 18562 15326
rect 18510 15250 18562 15262
rect 18734 15314 18786 15326
rect 18734 15250 18786 15262
rect 19182 15314 19234 15326
rect 20526 15314 20578 15326
rect 20290 15262 20302 15314
rect 20354 15262 20366 15314
rect 19182 15250 19234 15262
rect 20526 15250 20578 15262
rect 20750 15314 20802 15326
rect 20750 15250 20802 15262
rect 20974 15314 21026 15326
rect 24670 15314 24722 15326
rect 21298 15262 21310 15314
rect 21362 15262 21374 15314
rect 20974 15250 21026 15262
rect 24670 15250 24722 15262
rect 16718 15202 16770 15214
rect 14578 15150 14590 15202
rect 14642 15150 14654 15202
rect 16718 15138 16770 15150
rect 18062 15202 18114 15214
rect 18062 15138 18114 15150
rect 18622 15202 18674 15214
rect 24210 15150 24222 15202
rect 24274 15150 24286 15202
rect 18622 15138 18674 15150
rect 16270 15090 16322 15102
rect 17602 15038 17614 15090
rect 17666 15038 17678 15090
rect 16270 15026 16322 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 18734 14754 18786 14766
rect 18734 14690 18786 14702
rect 18958 14754 19010 14766
rect 18958 14690 19010 14702
rect 22990 14754 23042 14766
rect 22990 14690 23042 14702
rect 19182 14642 19234 14654
rect 15362 14590 15374 14642
rect 15426 14590 15438 14642
rect 17490 14590 17502 14642
rect 17554 14590 17566 14642
rect 19394 14590 19406 14642
rect 19458 14590 19470 14642
rect 19182 14578 19234 14590
rect 17950 14530 18002 14542
rect 14690 14478 14702 14530
rect 14754 14478 14766 14530
rect 17950 14466 18002 14478
rect 19406 14418 19458 14430
rect 18274 14366 18286 14418
rect 18338 14366 18350 14418
rect 19406 14354 19458 14366
rect 20526 14418 20578 14430
rect 20526 14354 20578 14366
rect 23102 14418 23154 14430
rect 23102 14354 23154 14366
rect 19630 14306 19682 14318
rect 19630 14242 19682 14254
rect 20414 14306 20466 14318
rect 20414 14242 20466 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 16382 13970 16434 13982
rect 16382 13906 16434 13918
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 24334 13970 24386 13982
rect 24334 13906 24386 13918
rect 40238 13858 40290 13870
rect 18162 13806 18174 13858
rect 18226 13806 18238 13858
rect 21746 13806 21758 13858
rect 21810 13806 21822 13858
rect 40238 13794 40290 13806
rect 17490 13694 17502 13746
rect 17554 13694 17566 13746
rect 21074 13694 21086 13746
rect 21138 13694 21150 13746
rect 20290 13582 20302 13634
rect 20354 13582 20366 13634
rect 23874 13582 23886 13634
rect 23938 13582 23950 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 17614 13074 17666 13086
rect 18610 13022 18622 13074
rect 18674 13022 18686 13074
rect 20738 13022 20750 13074
rect 20802 13022 20814 13074
rect 17614 13010 17666 13022
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 21310 12738 21362 12750
rect 21634 12686 21646 12738
rect 21698 12686 21710 12738
rect 21310 12674 21362 12686
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 26126 5234 26178 5246
rect 26126 5170 26178 5182
rect 25330 5070 25342 5122
rect 25394 5070 25406 5122
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 17714 4286 17726 4338
rect 17778 4286 17790 4338
rect 21074 4286 21086 4338
rect 21138 4286 21150 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 18734 4114 18786 4126
rect 18734 4050 18786 4062
rect 22094 4114 22146 4126
rect 22094 4050 22146 4062
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 22430 3666 22482 3678
rect 18162 3614 18174 3666
rect 18226 3614 18238 3666
rect 22430 3602 22482 3614
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 21410 3502 21422 3554
rect 21474 3502 21486 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18622 38222 18674 38274
rect 22094 38222 22146 38274
rect 25566 38222 25618 38274
rect 17950 37998 18002 38050
rect 21198 37998 21250 38050
rect 25006 37998 25058 38050
rect 27470 37886 27522 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18510 37438 18562 37490
rect 21422 37438 21474 37490
rect 26238 37438 26290 37490
rect 17614 37214 17666 37266
rect 20638 37214 20690 37266
rect 25230 37214 25282 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 18062 36654 18114 36706
rect 17390 36430 17442 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 17390 28702 17442 28754
rect 14590 28590 14642 28642
rect 18510 28590 18562 28642
rect 21758 28590 21810 28642
rect 15262 28478 15314 28530
rect 17726 28478 17778 28530
rect 18062 28478 18114 28530
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 15934 28030 15986 28082
rect 16718 28030 16770 28082
rect 17390 28030 17442 28082
rect 17726 28030 17778 28082
rect 16158 27918 16210 27970
rect 16270 27806 16322 27858
rect 16494 27806 16546 27858
rect 16830 27806 16882 27858
rect 18622 27806 18674 27858
rect 21758 27806 21810 27858
rect 19294 27694 19346 27746
rect 21422 27694 21474 27746
rect 22542 27694 22594 27746
rect 24670 27694 24722 27746
rect 25342 27694 25394 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 25454 27246 25506 27298
rect 20638 27134 20690 27186
rect 25118 27134 25170 27186
rect 40014 27134 40066 27186
rect 17838 27022 17890 27074
rect 22318 27022 22370 27074
rect 37662 27022 37714 27074
rect 18510 26910 18562 26962
rect 21422 26910 21474 26962
rect 21534 26910 21586 26962
rect 22990 26910 23042 26962
rect 25566 26910 25618 26962
rect 21198 26798 21250 26850
rect 26014 26798 26066 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17390 26462 17442 26514
rect 19070 26462 19122 26514
rect 19742 26462 19794 26514
rect 20526 26462 20578 26514
rect 21422 26462 21474 26514
rect 22654 26462 22706 26514
rect 23326 26462 23378 26514
rect 23438 26462 23490 26514
rect 23550 26462 23602 26514
rect 24334 26462 24386 26514
rect 24446 26462 24498 26514
rect 24558 26462 24610 26514
rect 18958 26350 19010 26402
rect 4286 26238 4338 26290
rect 15598 26238 15650 26290
rect 17726 26238 17778 26290
rect 19518 26238 19570 26290
rect 20190 26238 20242 26290
rect 20414 26238 20466 26290
rect 20638 26238 20690 26290
rect 21086 26238 21138 26290
rect 22542 26238 22594 26290
rect 23102 26238 23154 26290
rect 23214 26238 23266 26290
rect 24110 26238 24162 26290
rect 24222 26238 24274 26290
rect 25454 26238 25506 26290
rect 12686 26126 12738 26178
rect 14814 26126 14866 26178
rect 16046 26126 16098 26178
rect 16830 26126 16882 26178
rect 19630 26126 19682 26178
rect 26238 26126 26290 26178
rect 28366 26126 28418 26178
rect 1934 26014 1986 26066
rect 19182 26014 19234 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 2046 25566 2098 25618
rect 16382 25566 16434 25618
rect 16830 25566 16882 25618
rect 17502 25566 17554 25618
rect 26014 25566 26066 25618
rect 4286 25454 4338 25506
rect 13582 25454 13634 25506
rect 17054 25454 17106 25506
rect 26574 25454 26626 25506
rect 27022 25454 27074 25506
rect 27358 25454 27410 25506
rect 27806 25454 27858 25506
rect 14254 25342 14306 25394
rect 16718 25342 16770 25394
rect 27246 25342 27298 25394
rect 25118 25230 25170 25282
rect 25902 25230 25954 25282
rect 26126 25230 26178 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 14590 24894 14642 24946
rect 16158 24894 16210 24946
rect 17614 24894 17666 24946
rect 18398 24894 18450 24946
rect 22542 24894 22594 24946
rect 16270 24782 16322 24834
rect 18286 24782 18338 24834
rect 21310 24782 21362 24834
rect 22318 24782 22370 24834
rect 15934 24670 15986 24722
rect 17390 24670 17442 24722
rect 18062 24670 18114 24722
rect 18622 24670 18674 24722
rect 20750 24670 20802 24722
rect 21198 24670 21250 24722
rect 22206 24670 22258 24722
rect 37662 24670 37714 24722
rect 14702 24558 14754 24610
rect 17502 24558 17554 24610
rect 20974 24446 21026 24498
rect 40014 24446 40066 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 16270 24110 16322 24162
rect 16606 24110 16658 24162
rect 18958 24110 19010 24162
rect 28590 23998 28642 24050
rect 17614 23886 17666 23938
rect 25678 23886 25730 23938
rect 16830 23774 16882 23826
rect 17838 23774 17890 23826
rect 18622 23774 18674 23826
rect 18846 23774 18898 23826
rect 22542 23774 22594 23826
rect 23214 23774 23266 23826
rect 26462 23774 26514 23826
rect 22206 23662 22258 23714
rect 22430 23662 22482 23714
rect 22878 23662 22930 23714
rect 25342 23662 25394 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 16382 23326 16434 23378
rect 17726 23326 17778 23378
rect 18062 23326 18114 23378
rect 18846 23326 18898 23378
rect 19182 23326 19234 23378
rect 23774 23326 23826 23378
rect 26350 23326 26402 23378
rect 27358 23326 27410 23378
rect 27918 23326 27970 23378
rect 18622 23214 18674 23266
rect 19070 23214 19122 23266
rect 19630 23214 19682 23266
rect 23550 23214 23602 23266
rect 23998 23214 24050 23266
rect 27470 23214 27522 23266
rect 16046 23102 16098 23154
rect 19518 23102 19570 23154
rect 19854 23102 19906 23154
rect 20078 23102 20130 23154
rect 20414 23102 20466 23154
rect 21086 23102 21138 23154
rect 26238 23102 26290 23154
rect 26462 23102 26514 23154
rect 26910 23102 26962 23154
rect 27134 23102 27186 23154
rect 37662 23102 37714 23154
rect 15374 22990 15426 23042
rect 23214 22990 23266 23042
rect 24446 22990 24498 23042
rect 15486 22878 15538 22930
rect 23662 22878 23714 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 12910 22430 12962 22482
rect 13582 22430 13634 22482
rect 14030 22430 14082 22482
rect 27022 22430 27074 22482
rect 40014 22430 40066 22482
rect 10110 22318 10162 22370
rect 14590 22318 14642 22370
rect 15486 22318 15538 22370
rect 15934 22318 15986 22370
rect 16494 22318 16546 22370
rect 16830 22318 16882 22370
rect 17054 22318 17106 22370
rect 17726 22318 17778 22370
rect 21982 22318 22034 22370
rect 26798 22318 26850 22370
rect 37886 22318 37938 22370
rect 10782 22206 10834 22258
rect 25790 22206 25842 22258
rect 14142 22094 14194 22146
rect 14814 22094 14866 22146
rect 15598 22094 15650 22146
rect 16718 22094 16770 22146
rect 17390 22094 17442 22146
rect 17614 22094 17666 22146
rect 18846 22094 18898 22146
rect 19182 22094 19234 22146
rect 27134 22094 27186 22146
rect 27358 22094 27410 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14254 21758 14306 21810
rect 15038 21758 15090 21810
rect 17614 21758 17666 21810
rect 24110 21758 24162 21810
rect 11678 21646 11730 21698
rect 15374 21646 15426 21698
rect 15822 21646 15874 21698
rect 24334 21646 24386 21698
rect 11006 21534 11058 21586
rect 15710 21534 15762 21586
rect 15934 21534 15986 21586
rect 16270 21534 16322 21586
rect 17838 21534 17890 21586
rect 18174 21534 18226 21586
rect 23886 21534 23938 21586
rect 25790 21534 25842 21586
rect 37662 21534 37714 21586
rect 13806 21422 13858 21474
rect 20302 21422 20354 21474
rect 23998 21422 24050 21474
rect 25454 21422 25506 21474
rect 26574 21422 26626 21474
rect 28702 21422 28754 21474
rect 40014 21422 40066 21474
rect 17502 21310 17554 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 14702 20974 14754 21026
rect 14926 20974 14978 21026
rect 26798 20974 26850 21026
rect 14926 20862 14978 20914
rect 17950 20862 18002 20914
rect 23662 20862 23714 20914
rect 25790 20862 25842 20914
rect 27358 20862 27410 20914
rect 15486 20750 15538 20802
rect 15822 20750 15874 20802
rect 16158 20750 16210 20802
rect 18846 20750 18898 20802
rect 19630 20750 19682 20802
rect 19854 20750 19906 20802
rect 20190 20750 20242 20802
rect 21534 20750 21586 20802
rect 22206 20750 22258 20802
rect 22878 20750 22930 20802
rect 16718 20638 16770 20690
rect 18510 20638 18562 20690
rect 20078 20638 20130 20690
rect 21870 20638 21922 20690
rect 26238 20638 26290 20690
rect 26350 20638 26402 20690
rect 26686 20638 26738 20690
rect 26798 20638 26850 20690
rect 16046 20526 16098 20578
rect 16382 20526 16434 20578
rect 18174 20526 18226 20578
rect 19182 20526 19234 20578
rect 19966 20526 20018 20578
rect 22542 20526 22594 20578
rect 26014 20526 26066 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 15150 20190 15202 20242
rect 19070 20190 19122 20242
rect 19966 20190 20018 20242
rect 25902 20190 25954 20242
rect 15934 20078 15986 20130
rect 17726 20078 17778 20130
rect 18510 20078 18562 20130
rect 18622 20078 18674 20130
rect 19406 20078 19458 20130
rect 20526 20078 20578 20130
rect 20638 20078 20690 20130
rect 21534 20078 21586 20130
rect 21758 20078 21810 20130
rect 21982 20078 22034 20130
rect 22094 20078 22146 20130
rect 22318 20078 22370 20130
rect 24334 20078 24386 20130
rect 24670 20078 24722 20130
rect 25342 20078 25394 20130
rect 25790 20078 25842 20130
rect 26126 20078 26178 20130
rect 26350 20078 26402 20130
rect 26574 20078 26626 20130
rect 14814 19966 14866 20018
rect 15598 19966 15650 20018
rect 17390 19966 17442 20018
rect 18286 19966 18338 20018
rect 19294 19966 19346 20018
rect 19518 19966 19570 20018
rect 19742 19966 19794 20018
rect 20078 19966 20130 20018
rect 21422 19966 21474 20018
rect 25566 19966 25618 20018
rect 37662 19966 37714 20018
rect 13806 19854 13858 19906
rect 15038 19854 15090 19906
rect 16270 19854 16322 19906
rect 13918 19742 13970 19794
rect 20526 19742 20578 19794
rect 26238 19742 26290 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 15262 19294 15314 19346
rect 24782 19294 24834 19346
rect 28030 19294 28082 19346
rect 40014 19294 40066 19346
rect 13470 19182 13522 19234
rect 14478 19182 14530 19234
rect 14702 19182 14754 19234
rect 20078 19182 20130 19234
rect 21198 19182 21250 19234
rect 21422 19182 21474 19234
rect 21646 19182 21698 19234
rect 21870 19182 21922 19234
rect 22206 19182 22258 19234
rect 25230 19182 25282 19234
rect 37662 19182 37714 19234
rect 24334 19070 24386 19122
rect 24558 19070 24610 19122
rect 25902 19070 25954 19122
rect 13806 18958 13858 19010
rect 14254 18958 14306 19010
rect 14590 18958 14642 19010
rect 22542 18958 22594 19010
rect 23662 18958 23714 19010
rect 23998 18958 24050 19010
rect 24222 18958 24274 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 14814 18622 14866 18674
rect 19630 18622 19682 18674
rect 19966 18622 20018 18674
rect 21310 18622 21362 18674
rect 15038 18510 15090 18562
rect 15374 18510 15426 18562
rect 16830 18510 16882 18562
rect 17390 18510 17442 18562
rect 17726 18510 17778 18562
rect 18846 18510 18898 18562
rect 20638 18510 20690 18562
rect 20974 18510 21026 18562
rect 21086 18510 21138 18562
rect 4286 18398 4338 18450
rect 10670 18398 10722 18450
rect 14142 18398 14194 18450
rect 15262 18398 15314 18450
rect 16046 18398 16098 18450
rect 16606 18398 16658 18450
rect 18510 18398 18562 18450
rect 20302 18398 20354 18450
rect 25342 18398 25394 18450
rect 26014 18398 26066 18450
rect 11342 18286 11394 18338
rect 13470 18286 13522 18338
rect 13918 18286 13970 18338
rect 15038 18286 15090 18338
rect 16494 18286 16546 18338
rect 18174 18286 18226 18338
rect 24670 18286 24722 18338
rect 28142 18286 28194 18338
rect 1934 18174 1986 18226
rect 14478 18174 14530 18226
rect 16270 18174 16322 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 14366 17838 14418 17890
rect 14702 17838 14754 17890
rect 15598 17838 15650 17890
rect 16494 17838 16546 17890
rect 19182 17838 19234 17890
rect 13694 17726 13746 17778
rect 18958 17726 19010 17778
rect 15038 17614 15090 17666
rect 15262 17614 15314 17666
rect 15710 17614 15762 17666
rect 16158 17614 16210 17666
rect 16718 17614 16770 17666
rect 18622 17614 18674 17666
rect 19854 17614 19906 17666
rect 22318 17614 22370 17666
rect 14478 17502 14530 17554
rect 17390 17502 17442 17554
rect 20190 17502 20242 17554
rect 22766 17502 22818 17554
rect 15150 17390 15202 17442
rect 17054 17390 17106 17442
rect 18510 17390 18562 17442
rect 19518 17390 19570 17442
rect 22878 17390 22930 17442
rect 22990 17390 23042 17442
rect 23102 17390 23154 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 21198 17054 21250 17106
rect 21422 17054 21474 17106
rect 22542 17054 22594 17106
rect 23438 17054 23490 17106
rect 23662 17054 23714 17106
rect 13022 16942 13074 16994
rect 21534 16942 21586 16994
rect 21646 16942 21698 16994
rect 22654 16942 22706 16994
rect 23774 16942 23826 16994
rect 13694 16830 13746 16882
rect 14254 16830 14306 16882
rect 22318 16830 22370 16882
rect 22990 16830 23042 16882
rect 24222 16830 24274 16882
rect 10894 16718 10946 16770
rect 21982 16718 22034 16770
rect 22430 16718 22482 16770
rect 23550 16718 23602 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 18062 16270 18114 16322
rect 23998 16158 24050 16210
rect 26126 16158 26178 16210
rect 17278 16046 17330 16098
rect 17502 16046 17554 16098
rect 17726 16046 17778 16098
rect 19406 16046 19458 16098
rect 23214 16046 23266 16098
rect 19182 15934 19234 15986
rect 17614 15822 17666 15874
rect 18174 15822 18226 15874
rect 18286 15822 18338 15874
rect 26574 15822 26626 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 15038 15486 15090 15538
rect 21086 15486 21138 15538
rect 12462 15374 12514 15426
rect 17950 15374 18002 15426
rect 20078 15374 20130 15426
rect 22094 15374 22146 15426
rect 11790 15262 11842 15314
rect 16382 15262 16434 15314
rect 16606 15262 16658 15314
rect 17614 15262 17666 15314
rect 18174 15262 18226 15314
rect 18510 15262 18562 15314
rect 18734 15262 18786 15314
rect 19182 15262 19234 15314
rect 20302 15262 20354 15314
rect 20526 15262 20578 15314
rect 20750 15262 20802 15314
rect 20974 15262 21026 15314
rect 21310 15262 21362 15314
rect 24670 15262 24722 15314
rect 14590 15150 14642 15202
rect 16718 15150 16770 15202
rect 18062 15150 18114 15202
rect 18622 15150 18674 15202
rect 24222 15150 24274 15202
rect 16270 15038 16322 15090
rect 17614 15038 17666 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 18734 14702 18786 14754
rect 18958 14702 19010 14754
rect 22990 14702 23042 14754
rect 15374 14590 15426 14642
rect 17502 14590 17554 14642
rect 19182 14590 19234 14642
rect 19406 14590 19458 14642
rect 14702 14478 14754 14530
rect 17950 14478 18002 14530
rect 18286 14366 18338 14418
rect 19406 14366 19458 14418
rect 20526 14366 20578 14418
rect 23102 14366 23154 14418
rect 19630 14254 19682 14306
rect 20414 14254 20466 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 16382 13918 16434 13970
rect 16830 13918 16882 13970
rect 24334 13918 24386 13970
rect 18174 13806 18226 13858
rect 21758 13806 21810 13858
rect 40238 13806 40290 13858
rect 17502 13694 17554 13746
rect 21086 13694 21138 13746
rect 20302 13582 20354 13634
rect 23886 13582 23938 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17614 13022 17666 13074
rect 18622 13022 18674 13074
rect 20750 13022 20802 13074
rect 17838 12910 17890 12962
rect 21310 12686 21362 12738
rect 21646 12686 21698 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 26126 5182 26178 5234
rect 25342 5070 25394 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 17726 4286 17778 4338
rect 21086 4286 21138 4338
rect 25230 4286 25282 4338
rect 18734 4062 18786 4114
rect 22094 4062 22146 4114
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18174 3614 18226 3666
rect 22430 3614 22482 3666
rect 25566 3614 25618 3666
rect 19742 3502 19794 3554
rect 21422 3502 21474 3554
rect 24558 3502 24610 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 16800 41200 16912 42000
rect 17472 41200 17584 42000
rect 18144 41200 18256 42000
rect 20160 41200 20272 42000
rect 20832 41200 20944 42000
rect 24192 41200 24304 42000
rect 24864 41200 24976 42000
rect 26208 41200 26320 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 16828 36708 16884 41200
rect 17500 37492 17556 41200
rect 18172 38276 18228 41200
rect 18620 38276 18676 38286
rect 18172 38274 18676 38276
rect 18172 38222 18622 38274
rect 18674 38222 18676 38274
rect 18172 38220 18676 38222
rect 18620 38210 18676 38220
rect 17500 37426 17556 37436
rect 17948 38050 18004 38062
rect 17948 37998 17950 38050
rect 18002 37998 18004 38050
rect 16828 36642 16884 36652
rect 17612 37266 17668 37278
rect 17612 37214 17614 37266
rect 17666 37214 17668 37266
rect 17388 36482 17444 36494
rect 17388 36430 17390 36482
rect 17442 36430 17444 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 17388 28754 17444 36430
rect 17388 28702 17390 28754
rect 17442 28702 17444 28754
rect 14588 28644 14644 28654
rect 14588 28550 14644 28588
rect 15260 28532 15316 28542
rect 16716 28532 16772 28542
rect 15260 28530 15988 28532
rect 15260 28478 15262 28530
rect 15314 28478 15988 28530
rect 15260 28476 15988 28478
rect 15260 28466 15316 28476
rect 4172 28308 4228 28318
rect 1932 26066 1988 26078
rect 1932 26014 1934 26066
rect 1986 26014 1988 26066
rect 1932 25620 1988 26014
rect 1932 25554 1988 25564
rect 2044 25618 2100 25630
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 24948 2100 25566
rect 2044 24882 2100 24892
rect 4172 20580 4228 28252
rect 15932 28082 15988 28476
rect 15932 28030 15934 28082
rect 15986 28030 15988 28082
rect 15932 28018 15988 28030
rect 16716 28082 16772 28476
rect 16716 28030 16718 28082
rect 16770 28030 16772 28082
rect 16716 28018 16772 28030
rect 17388 28532 17444 28702
rect 17388 28082 17444 28476
rect 17388 28030 17390 28082
rect 17442 28030 17444 28082
rect 17388 28018 17444 28030
rect 17500 28644 17556 28654
rect 16156 27972 16212 27982
rect 16044 27970 16212 27972
rect 16044 27918 16158 27970
rect 16210 27918 16212 27970
rect 16044 27916 16212 27918
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 16044 26908 16100 27916
rect 16156 27906 16212 27916
rect 16268 27860 16324 27870
rect 16492 27860 16548 27870
rect 16268 27858 16548 27860
rect 16268 27806 16270 27858
rect 16322 27806 16494 27858
rect 16546 27806 16548 27858
rect 16268 27804 16548 27806
rect 16268 27794 16324 27804
rect 16492 27794 16548 27804
rect 16828 27858 16884 27870
rect 16828 27806 16830 27858
rect 16882 27806 16884 27858
rect 16828 26964 16884 27806
rect 16044 26852 16212 26908
rect 16828 26898 16884 26908
rect 17388 26964 17444 26974
rect 4284 26292 4340 26302
rect 4284 26198 4340 26236
rect 12684 26292 12740 26302
rect 12684 26178 12740 26236
rect 15596 26290 15652 26302
rect 15596 26238 15598 26290
rect 15650 26238 15652 26290
rect 12684 26126 12686 26178
rect 12738 26126 12740 26178
rect 12684 26114 12740 26126
rect 13580 26180 13636 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4284 25506 4340 25518
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 25396 4340 25454
rect 4284 25330 4340 25340
rect 13580 25506 13636 26124
rect 14812 26178 14868 26190
rect 14812 26126 14814 26178
rect 14866 26126 14868 26178
rect 14812 25732 14868 26126
rect 15596 26180 15652 26238
rect 15596 26114 15652 26124
rect 15932 26292 15988 26302
rect 14812 25666 14868 25676
rect 15260 26068 15316 26078
rect 13580 25454 13582 25506
rect 13634 25454 13636 25506
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 12908 22484 12964 22494
rect 12908 22390 12964 22428
rect 13580 22482 13636 25454
rect 14252 25396 14308 25406
rect 14252 25394 14644 25396
rect 14252 25342 14254 25394
rect 14306 25342 14644 25394
rect 14252 25340 14644 25342
rect 14252 25330 14308 25340
rect 14588 24946 14644 25340
rect 14588 24894 14590 24946
rect 14642 24894 14644 24946
rect 14588 24882 14644 24894
rect 14700 24610 14756 24622
rect 14700 24558 14702 24610
rect 14754 24558 14756 24610
rect 14700 24164 14756 24558
rect 14700 24098 14756 24108
rect 13580 22430 13582 22482
rect 13634 22430 13636 22482
rect 10108 22370 10164 22382
rect 10108 22318 10110 22370
rect 10162 22318 10164 22370
rect 10108 21812 10164 22318
rect 10108 21746 10164 21756
rect 10780 22258 10836 22270
rect 10780 22206 10782 22258
rect 10834 22206 10836 22258
rect 10780 21700 10836 22206
rect 11676 21924 11732 21934
rect 10780 21634 10836 21644
rect 11004 21812 11060 21822
rect 11004 21588 11060 21756
rect 11676 21698 11732 21868
rect 11676 21646 11678 21698
rect 11730 21646 11732 21698
rect 11676 21634 11732 21646
rect 13580 21812 13636 22430
rect 14028 22484 14084 22494
rect 14028 22390 14084 22428
rect 14588 22484 14644 22494
rect 14588 22370 14644 22428
rect 14588 22318 14590 22370
rect 14642 22318 14644 22370
rect 14588 22306 14644 22318
rect 14924 22484 14980 22494
rect 14140 22148 14196 22158
rect 14140 22054 14196 22092
rect 14812 22146 14868 22158
rect 14812 22094 14814 22146
rect 14866 22094 14868 22146
rect 10892 21586 11060 21588
rect 10892 21534 11006 21586
rect 11058 21534 11060 21586
rect 10892 21532 11060 21534
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4172 20514 4228 20524
rect 10892 20188 10948 21532
rect 11004 21522 11060 21532
rect 13580 20356 13636 21756
rect 14252 21812 14308 21822
rect 14252 21718 14308 21756
rect 13580 20188 13636 20300
rect 10668 20132 10948 20188
rect 13356 20132 13636 20188
rect 13804 21474 13860 21486
rect 13804 21422 13806 21474
rect 13858 21422 13860 21474
rect 13804 20188 13860 21422
rect 14700 21028 14756 21038
rect 14476 21026 14756 21028
rect 14476 20974 14702 21026
rect 14754 20974 14756 21026
rect 14476 20972 14756 20974
rect 13804 20132 13972 20188
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4284 18450 4340 18462
rect 4284 18398 4286 18450
rect 4338 18398 4340 18450
rect 1932 18228 1988 18238
rect 1932 18134 1988 18172
rect 4284 17668 4340 18398
rect 10668 18450 10724 20132
rect 10668 18398 10670 18450
rect 10722 18398 10724 18450
rect 10668 18386 10724 18398
rect 11340 18340 11396 18350
rect 11340 18246 11396 18284
rect 13356 18116 13412 20132
rect 13916 20020 13972 20132
rect 13916 19954 13972 19964
rect 13804 19906 13860 19918
rect 13804 19854 13806 19906
rect 13858 19854 13860 19906
rect 13804 19348 13860 19854
rect 13916 19794 13972 19806
rect 13916 19742 13918 19794
rect 13970 19742 13972 19794
rect 13916 19460 13972 19742
rect 13916 19394 13972 19404
rect 13468 19292 13860 19348
rect 13468 19234 13524 19292
rect 13468 19182 13470 19234
rect 13522 19182 13524 19234
rect 13468 18338 13524 19182
rect 14476 19234 14532 20972
rect 14700 20962 14756 20972
rect 14812 21028 14868 22094
rect 14812 20018 14868 20972
rect 14924 21026 14980 22428
rect 15260 22484 15316 26012
rect 15932 24722 15988 26236
rect 16044 26180 16100 26190
rect 16044 26086 16100 26124
rect 16156 25508 16212 26852
rect 17388 26514 17444 26908
rect 17388 26462 17390 26514
rect 17442 26462 17444 26514
rect 17388 26450 17444 26462
rect 16828 26178 16884 26190
rect 16828 26126 16830 26178
rect 16882 26126 16884 26178
rect 16828 26068 16884 26126
rect 16828 26002 16884 26012
rect 17500 26180 17556 28588
rect 17612 28084 17668 37214
rect 17948 31948 18004 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18508 37492 18564 37502
rect 18508 37398 18564 37436
rect 20188 37492 20244 41200
rect 20860 38276 20916 41200
rect 20860 38210 20916 38220
rect 22092 38276 22148 38286
rect 22092 38182 22148 38220
rect 24220 38276 24276 41200
rect 24220 38210 24276 38220
rect 20188 37426 20244 37436
rect 21196 38050 21252 38062
rect 21196 37998 21198 38050
rect 21250 37998 21252 38050
rect 20636 37266 20692 37278
rect 20636 37214 20638 37266
rect 20690 37214 20692 37266
rect 18060 36708 18116 36718
rect 18060 36614 18116 36652
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 17948 31892 18116 31948
rect 17724 28532 17780 28542
rect 17724 28438 17780 28476
rect 18060 28530 18116 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 18508 28644 18564 28654
rect 18508 28550 18564 28588
rect 18060 28478 18062 28530
rect 18114 28478 18116 28530
rect 18060 28466 18116 28478
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 17724 28084 17780 28094
rect 17612 28082 17780 28084
rect 17612 28030 17726 28082
rect 17778 28030 17780 28082
rect 17612 28028 17780 28030
rect 17724 28018 17780 28028
rect 17836 27860 17892 27870
rect 17836 27074 17892 27804
rect 18620 27860 18676 27870
rect 18620 27766 18676 27804
rect 17836 27022 17838 27074
rect 17890 27022 17892 27074
rect 17836 27010 17892 27022
rect 19292 27746 19348 27758
rect 19292 27694 19294 27746
rect 19346 27694 19348 27746
rect 18508 26964 18564 26974
rect 18508 26962 18900 26964
rect 18508 26910 18510 26962
rect 18562 26910 18900 26962
rect 18508 26908 18900 26910
rect 18508 26898 18564 26908
rect 18844 26852 19124 26908
rect 19068 26514 19124 26852
rect 19292 26852 19348 27694
rect 20636 27186 20692 37214
rect 21196 31948 21252 37998
rect 21420 37492 21476 37502
rect 21420 37398 21476 37436
rect 24892 37492 24948 41200
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 25004 38052 25060 38062
rect 25004 38050 25172 38052
rect 25004 37998 25006 38050
rect 25058 37998 25172 38050
rect 25004 37996 25172 37998
rect 25004 37986 25060 37996
rect 24892 37426 24948 37436
rect 21196 31892 21476 31948
rect 20636 27134 20638 27186
rect 20690 27134 20692 27186
rect 19292 26786 19348 26796
rect 20524 26852 20580 26862
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19068 26462 19070 26514
rect 19122 26462 19124 26514
rect 19068 26450 19124 26462
rect 19740 26516 19796 26526
rect 19740 26422 19796 26460
rect 20524 26514 20580 26796
rect 20524 26462 20526 26514
rect 20578 26462 20580 26514
rect 20524 26450 20580 26462
rect 20636 26516 20692 27134
rect 21308 27860 21364 27870
rect 20636 26450 20692 26460
rect 21196 26850 21252 26862
rect 21196 26798 21198 26850
rect 21250 26798 21252 26850
rect 18956 26402 19012 26414
rect 18956 26350 18958 26402
rect 19010 26350 19012 26402
rect 16380 25732 16436 25742
rect 16380 25618 16436 25676
rect 16380 25566 16382 25618
rect 16434 25566 16436 25618
rect 16380 25554 16436 25566
rect 16828 25620 16884 25630
rect 16828 25526 16884 25564
rect 17500 25618 17556 26124
rect 17724 26290 17780 26302
rect 17724 26238 17726 26290
rect 17778 26238 17780 26290
rect 17724 26068 17780 26238
rect 17724 26002 17780 26012
rect 17500 25566 17502 25618
rect 17554 25566 17556 25618
rect 17500 25554 17556 25566
rect 17612 25732 17668 25742
rect 15932 24670 15934 24722
rect 15986 24670 15988 24722
rect 15932 24658 15988 24670
rect 16044 25452 16212 25508
rect 17052 25508 17108 25518
rect 17052 25506 17220 25508
rect 17052 25454 17054 25506
rect 17106 25454 17220 25506
rect 17052 25452 17220 25454
rect 16044 25060 16100 25452
rect 17052 25442 17108 25452
rect 16716 25396 16772 25406
rect 16044 23548 16100 25004
rect 16156 25394 16772 25396
rect 16156 25342 16718 25394
rect 16770 25342 16772 25394
rect 16156 25340 16772 25342
rect 16156 24946 16212 25340
rect 16716 25330 16772 25340
rect 16156 24894 16158 24946
rect 16210 24894 16212 24946
rect 16156 24882 16212 24894
rect 16268 24948 16324 24958
rect 16268 24834 16324 24892
rect 16268 24782 16270 24834
rect 16322 24782 16324 24834
rect 16268 24770 16324 24782
rect 16604 24612 16660 24622
rect 16268 24164 16324 24174
rect 16268 24070 16324 24108
rect 16604 24162 16660 24556
rect 16604 24110 16606 24162
rect 16658 24110 16660 24162
rect 16604 24098 16660 24110
rect 16828 23828 16884 23838
rect 16828 23826 17108 23828
rect 16828 23774 16830 23826
rect 16882 23774 17108 23826
rect 16828 23772 17108 23774
rect 16828 23762 16884 23772
rect 17052 23548 17108 23772
rect 16044 23492 16324 23548
rect 16044 23154 16100 23166
rect 16044 23102 16046 23154
rect 16098 23102 16100 23154
rect 15260 22418 15316 22428
rect 15372 23042 15428 23054
rect 15372 22990 15374 23042
rect 15426 22990 15428 23042
rect 15036 22148 15092 22158
rect 15036 21810 15092 22092
rect 15372 21924 15428 22990
rect 15484 22932 15540 22942
rect 16044 22932 16100 23102
rect 15484 22930 16100 22932
rect 15484 22878 15486 22930
rect 15538 22878 16100 22930
rect 15484 22876 16100 22878
rect 15484 22370 15540 22876
rect 15484 22318 15486 22370
rect 15538 22318 15540 22370
rect 15484 22306 15540 22318
rect 15596 22484 15652 22494
rect 15596 22146 15652 22428
rect 15932 22372 15988 22382
rect 15932 22370 16100 22372
rect 15932 22318 15934 22370
rect 15986 22318 16100 22370
rect 15932 22316 16100 22318
rect 15932 22306 15988 22316
rect 15596 22094 15598 22146
rect 15650 22094 15652 22146
rect 15596 22082 15652 22094
rect 16044 22148 16100 22316
rect 15036 21758 15038 21810
rect 15090 21758 15092 21810
rect 15036 21746 15092 21758
rect 15260 21868 15428 21924
rect 14924 20974 14926 21026
rect 14978 20974 14980 21026
rect 14924 20914 14980 20974
rect 14924 20862 14926 20914
rect 14978 20862 14980 20914
rect 14924 20850 14980 20862
rect 15260 20804 15316 21868
rect 15372 21698 15428 21710
rect 15372 21646 15374 21698
rect 15426 21646 15428 21698
rect 15372 21140 15428 21646
rect 15820 21700 15876 21710
rect 15820 21606 15876 21644
rect 15708 21586 15764 21598
rect 15708 21534 15710 21586
rect 15762 21534 15764 21586
rect 15708 21364 15764 21534
rect 15708 21298 15764 21308
rect 15932 21586 15988 21598
rect 15932 21534 15934 21586
rect 15986 21534 15988 21586
rect 15932 21140 15988 21534
rect 15372 21084 15988 21140
rect 15484 20804 15540 20814
rect 15260 20802 15540 20804
rect 15260 20750 15486 20802
rect 15538 20750 15540 20802
rect 15260 20748 15540 20750
rect 15148 20242 15204 20254
rect 15148 20190 15150 20242
rect 15202 20190 15204 20242
rect 15148 20132 15204 20190
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14812 19954 14868 19966
rect 15036 20020 15092 20030
rect 15036 19906 15092 19964
rect 15036 19854 15038 19906
rect 15090 19854 15092 19906
rect 15036 19842 15092 19854
rect 15148 19348 15204 20076
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14476 19170 14532 19182
rect 14700 19292 15204 19348
rect 15260 20244 15316 20254
rect 15260 19346 15316 20188
rect 15372 20020 15428 20748
rect 15484 20738 15540 20748
rect 15708 20580 15764 21084
rect 15820 20804 15876 20814
rect 16044 20804 16100 22092
rect 16268 21586 16324 23492
rect 16940 23492 17108 23548
rect 17164 23548 17220 25452
rect 17612 24946 17668 25676
rect 18284 25060 18340 25070
rect 17612 24894 17614 24946
rect 17666 24894 17668 24946
rect 17612 24882 17668 24894
rect 17836 24948 17892 24958
rect 17388 24722 17444 24734
rect 17388 24670 17390 24722
rect 17442 24670 17444 24722
rect 17388 23716 17444 24670
rect 17500 24612 17556 24622
rect 17500 24518 17556 24556
rect 17388 23650 17444 23660
rect 17612 23938 17668 23950
rect 17612 23886 17614 23938
rect 17666 23886 17668 23938
rect 17612 23828 17668 23886
rect 16380 23380 16436 23390
rect 16380 23286 16436 23324
rect 16268 21534 16270 21586
rect 16322 21534 16324 21586
rect 15820 20802 16100 20804
rect 15820 20750 15822 20802
rect 15874 20750 16100 20802
rect 15820 20748 16100 20750
rect 16156 20804 16212 20814
rect 15820 20738 15876 20748
rect 16156 20710 16212 20748
rect 15708 20524 15876 20580
rect 15372 19954 15428 19964
rect 15596 20132 15652 20142
rect 15596 20018 15652 20076
rect 15596 19966 15598 20018
rect 15650 19966 15652 20018
rect 15596 19954 15652 19966
rect 15820 19908 15876 20524
rect 16044 20578 16100 20590
rect 16044 20526 16046 20578
rect 16098 20526 16100 20578
rect 15820 19842 15876 19852
rect 15932 20132 15988 20142
rect 15260 19294 15262 19346
rect 15314 19294 15316 19346
rect 14700 19234 14756 19292
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14700 19170 14756 19182
rect 13468 18286 13470 18338
rect 13522 18286 13524 18338
rect 13468 18274 13524 18286
rect 13804 19010 13860 19022
rect 13804 18958 13806 19010
rect 13858 18958 13860 19010
rect 13804 18228 13860 18958
rect 14252 19010 14308 19022
rect 14252 18958 14254 19010
rect 14306 18958 14308 19010
rect 14140 18676 14196 18686
rect 14140 18450 14196 18620
rect 14140 18398 14142 18450
rect 14194 18398 14196 18450
rect 14140 18386 14196 18398
rect 14252 18452 14308 18958
rect 13916 18340 13972 18350
rect 13916 18246 13972 18284
rect 13804 18162 13860 18172
rect 4476 18060 4740 18070
rect 13356 18060 13748 18116
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 13692 17778 13748 18060
rect 13692 17726 13694 17778
rect 13746 17726 13748 17778
rect 4284 17602 4340 17612
rect 10892 17668 10948 17678
rect 10892 16770 10948 17612
rect 13020 17444 13076 17454
rect 13020 16994 13076 17388
rect 13020 16942 13022 16994
rect 13074 16942 13076 16994
rect 13020 16930 13076 16942
rect 13692 16884 13748 17726
rect 14252 17668 14308 18396
rect 14588 19010 14644 19022
rect 14588 18958 14590 19010
rect 14642 18958 14644 19010
rect 14364 18340 14420 18350
rect 14364 17890 14420 18284
rect 14364 17838 14366 17890
rect 14418 17838 14420 17890
rect 14364 17826 14420 17838
rect 14476 18226 14532 18238
rect 14476 18174 14478 18226
rect 14530 18174 14532 18226
rect 14476 17780 14532 18174
rect 14476 17714 14532 17724
rect 14252 17602 14308 17612
rect 14588 17668 14644 18958
rect 14812 18676 14868 19292
rect 15260 19282 15316 19294
rect 14812 18582 14868 18620
rect 15036 18564 15092 18574
rect 14924 18562 15092 18564
rect 14924 18510 15038 18562
rect 15090 18510 15092 18562
rect 14924 18508 15092 18510
rect 14924 18452 14980 18508
rect 15036 18498 15092 18508
rect 15372 18564 15428 18574
rect 15372 18470 15428 18508
rect 14924 18386 14980 18396
rect 15260 18450 15316 18462
rect 15260 18398 15262 18450
rect 15314 18398 15316 18450
rect 14700 18340 14756 18350
rect 14700 17890 14756 18284
rect 14700 17838 14702 17890
rect 14754 17838 14756 17890
rect 14700 17826 14756 17838
rect 15036 18338 15092 18350
rect 15036 18286 15038 18338
rect 15090 18286 15092 18338
rect 14588 17602 14644 17612
rect 15036 17666 15092 18286
rect 15260 18340 15316 18398
rect 15260 18274 15316 18284
rect 15932 18004 15988 20076
rect 16044 19460 16100 20526
rect 16268 19906 16324 21534
rect 16492 22370 16548 22382
rect 16492 22318 16494 22370
rect 16546 22318 16548 22370
rect 16492 22148 16548 22318
rect 16828 22370 16884 22382
rect 16828 22318 16830 22370
rect 16882 22318 16884 22370
rect 16380 20578 16436 20590
rect 16380 20526 16382 20578
rect 16434 20526 16436 20578
rect 16380 20132 16436 20526
rect 16380 20066 16436 20076
rect 16268 19854 16270 19906
rect 16322 19854 16324 19906
rect 16268 19684 16324 19854
rect 16268 19618 16324 19628
rect 16492 19460 16548 22092
rect 16716 22146 16772 22158
rect 16716 22094 16718 22146
rect 16770 22094 16772 22146
rect 16716 21924 16772 22094
rect 16716 21858 16772 21868
rect 16716 21364 16772 21374
rect 16828 21364 16884 22318
rect 16940 22372 16996 23492
rect 17164 23482 17220 23492
rect 17612 23380 17668 23772
rect 17836 23826 17892 24892
rect 18284 24834 18340 25004
rect 18956 25060 19012 26350
rect 19516 26292 19572 26302
rect 18956 24994 19012 25004
rect 19068 26290 19572 26292
rect 19068 26238 19518 26290
rect 19570 26238 19572 26290
rect 19068 26236 19572 26238
rect 18396 24948 18452 24958
rect 18396 24854 18452 24892
rect 19068 24948 19124 26236
rect 19516 26226 19572 26236
rect 20188 26292 20244 26302
rect 20188 26198 20244 26236
rect 20412 26290 20468 26302
rect 20412 26238 20414 26290
rect 20466 26238 20468 26290
rect 19628 26178 19684 26190
rect 19628 26126 19630 26178
rect 19682 26126 19684 26178
rect 19180 26068 19236 26078
rect 19628 26068 19684 26126
rect 19180 26066 19684 26068
rect 19180 26014 19182 26066
rect 19234 26014 19684 26066
rect 19180 26012 19684 26014
rect 19180 26002 19236 26012
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19068 24882 19124 24892
rect 18284 24782 18286 24834
rect 18338 24782 18340 24834
rect 18284 24770 18340 24782
rect 18732 24836 18788 24846
rect 18060 24724 18116 24734
rect 18620 24724 18676 24734
rect 17836 23774 17838 23826
rect 17890 23774 17892 23826
rect 17836 23604 17892 23774
rect 17836 23538 17892 23548
rect 17948 24668 18060 24724
rect 17724 23380 17780 23390
rect 17668 23378 17780 23380
rect 17668 23326 17726 23378
rect 17778 23326 17780 23378
rect 17668 23324 17780 23326
rect 17612 23286 17668 23324
rect 17052 22372 17108 22382
rect 16940 22370 17556 22372
rect 16940 22318 17054 22370
rect 17106 22318 17556 22370
rect 16940 22316 17556 22318
rect 17052 22306 17108 22316
rect 17388 22148 17444 22158
rect 17388 22054 17444 22092
rect 17500 21812 17556 22316
rect 17724 22370 17780 23324
rect 17724 22318 17726 22370
rect 17778 22318 17780 22370
rect 17724 22306 17780 22318
rect 17948 22260 18004 24668
rect 18060 24630 18116 24668
rect 18508 24722 18676 24724
rect 18508 24670 18622 24722
rect 18674 24670 18676 24722
rect 18508 24668 18676 24670
rect 17836 22204 18004 22260
rect 18060 23716 18116 23726
rect 18060 23378 18116 23660
rect 18060 23326 18062 23378
rect 18114 23326 18116 23378
rect 17612 22148 17668 22158
rect 17836 22148 17892 22204
rect 17612 22146 17892 22148
rect 17612 22094 17614 22146
rect 17666 22094 17892 22146
rect 17612 22092 17892 22094
rect 17612 22082 17668 22092
rect 17612 21812 17668 21822
rect 17500 21810 17668 21812
rect 17500 21758 17614 21810
rect 17666 21758 17668 21810
rect 17500 21756 17668 21758
rect 17612 21746 17668 21756
rect 18060 21812 18116 23326
rect 18508 23380 18564 24668
rect 18620 24658 18676 24668
rect 18620 23828 18676 23838
rect 18620 23734 18676 23772
rect 18508 23314 18564 23324
rect 18620 23604 18676 23614
rect 18620 23266 18676 23548
rect 18620 23214 18622 23266
rect 18674 23214 18676 23266
rect 18620 23202 18676 23214
rect 18732 23380 18788 24780
rect 18844 24724 18900 24734
rect 18844 23828 18900 24668
rect 18956 24612 19012 24622
rect 18956 24162 19012 24556
rect 19740 24164 19796 24174
rect 18956 24110 18958 24162
rect 19010 24110 19012 24162
rect 18956 24098 19012 24110
rect 19628 24108 19740 24164
rect 18844 23826 19012 23828
rect 18844 23774 18846 23826
rect 18898 23774 19012 23826
rect 18844 23772 19012 23774
rect 18844 23762 18900 23772
rect 18844 23380 18900 23390
rect 18732 23378 18900 23380
rect 18732 23326 18846 23378
rect 18898 23326 18900 23378
rect 18732 23324 18900 23326
rect 18060 21746 18116 21756
rect 17836 21588 17892 21598
rect 18172 21588 18228 21598
rect 17836 21494 17892 21532
rect 17948 21586 18228 21588
rect 17948 21534 18174 21586
rect 18226 21534 18228 21586
rect 17948 21532 18228 21534
rect 16772 21308 16884 21364
rect 17500 21364 17556 21374
rect 16716 20690 16772 21308
rect 17500 21270 17556 21308
rect 16716 20638 16718 20690
rect 16770 20638 16772 20690
rect 16716 20626 16772 20638
rect 17948 20914 18004 21532
rect 18172 21522 18228 21532
rect 17948 20862 17950 20914
rect 18002 20862 18004 20914
rect 17948 20580 18004 20862
rect 18508 20692 18564 20702
rect 18732 20692 18788 23324
rect 18844 23314 18900 23324
rect 18508 20690 18732 20692
rect 18508 20638 18510 20690
rect 18562 20638 18732 20690
rect 18508 20636 18732 20638
rect 18508 20626 18564 20636
rect 18732 20598 18788 20636
rect 18844 22146 18900 22158
rect 18844 22094 18846 22146
rect 18898 22094 18900 22146
rect 18844 21028 18900 22094
rect 18844 20802 18900 20972
rect 18844 20750 18846 20802
rect 18898 20750 18900 20802
rect 17948 20514 18004 20524
rect 18172 20578 18228 20590
rect 18172 20526 18174 20578
rect 18226 20526 18228 20578
rect 17724 20132 17780 20142
rect 17724 20038 17780 20076
rect 17388 20020 17444 20030
rect 17388 19926 17444 19964
rect 16044 19394 16100 19404
rect 16156 19404 16548 19460
rect 16828 19684 16884 19694
rect 16044 18452 16100 18462
rect 16156 18452 16212 19404
rect 16828 18562 16884 19628
rect 17388 19460 17444 19470
rect 16828 18510 16830 18562
rect 16882 18510 16884 18562
rect 16828 18498 16884 18510
rect 17276 18564 17332 18574
rect 16044 18450 16212 18452
rect 16044 18398 16046 18450
rect 16098 18398 16212 18450
rect 16044 18396 16212 18398
rect 16604 18450 16660 18462
rect 16604 18398 16606 18450
rect 16658 18398 16660 18450
rect 16044 18386 16100 18396
rect 16492 18340 16548 18350
rect 16380 18338 16548 18340
rect 16380 18286 16494 18338
rect 16546 18286 16548 18338
rect 16380 18284 16548 18286
rect 16268 18228 16324 18238
rect 16268 18134 16324 18172
rect 15932 17948 16212 18004
rect 15596 17890 15652 17902
rect 15596 17838 15598 17890
rect 15650 17838 15652 17890
rect 15036 17614 15038 17666
rect 15090 17614 15092 17666
rect 15036 17602 15092 17614
rect 15260 17668 15316 17678
rect 15260 17574 15316 17612
rect 14476 17556 14532 17566
rect 14476 17462 14532 17500
rect 15148 17444 15204 17454
rect 15596 17444 15652 17838
rect 15708 17668 15764 17678
rect 15708 17574 15764 17612
rect 16156 17668 16212 17948
rect 16156 17574 16212 17612
rect 16380 17444 16436 18284
rect 16492 18274 16548 18284
rect 16492 18116 16548 18126
rect 16492 17890 16548 18060
rect 16492 17838 16494 17890
rect 16546 17838 16548 17890
rect 16492 17826 16548 17838
rect 16604 17668 16660 18398
rect 17276 17780 17332 18508
rect 17388 18562 17444 19404
rect 18060 19012 18116 19022
rect 17388 18510 17390 18562
rect 17442 18510 17444 18562
rect 17388 18498 17444 18510
rect 17724 18564 17780 18574
rect 17276 17714 17332 17724
rect 16604 17602 16660 17612
rect 16716 17666 16772 17678
rect 16716 17614 16718 17666
rect 16770 17614 16772 17666
rect 15596 17388 16436 17444
rect 15148 17350 15204 17388
rect 14252 16884 14308 16894
rect 13692 16882 14308 16884
rect 13692 16830 13694 16882
rect 13746 16830 14254 16882
rect 14306 16830 14308 16882
rect 13692 16828 14308 16830
rect 13692 16818 13748 16828
rect 10892 16718 10894 16770
rect 10946 16718 10948 16770
rect 10892 16706 10948 16718
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 12460 16100 12516 16110
rect 11788 15540 11844 15550
rect 11788 15314 11844 15484
rect 12460 15426 12516 16044
rect 14252 15540 14308 16828
rect 14252 15474 14308 15484
rect 14588 16884 14644 16894
rect 12460 15374 12462 15426
rect 12514 15374 12516 15426
rect 12460 15362 12516 15374
rect 11788 15262 11790 15314
rect 11842 15262 11844 15314
rect 11788 15250 11844 15262
rect 14588 15202 14644 16828
rect 14588 15150 14590 15202
rect 14642 15150 14644 15202
rect 14588 15138 14644 15150
rect 14700 15540 14756 15550
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 14700 14532 14756 15484
rect 15036 15540 15092 15550
rect 15036 15446 15092 15484
rect 16380 15314 16436 17388
rect 16716 17444 16772 17614
rect 17388 17668 17444 17678
rect 17724 17668 17780 18508
rect 17388 17554 17444 17612
rect 17388 17502 17390 17554
rect 17442 17502 17444 17554
rect 17388 17490 17444 17502
rect 17500 17612 17780 17668
rect 17836 17780 17892 17790
rect 17052 17444 17108 17454
rect 16716 17442 17108 17444
rect 16716 17390 17054 17442
rect 17106 17390 17108 17442
rect 16716 17388 17108 17390
rect 16716 16884 16772 17388
rect 17052 17378 17108 17388
rect 16716 16818 16772 16828
rect 17276 16098 17332 16110
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 17276 15876 17332 16046
rect 17500 16100 17556 17612
rect 17500 16006 17556 16044
rect 17724 16100 17780 16110
rect 17836 16100 17892 17724
rect 18060 16324 18116 18956
rect 18172 18338 18228 20526
rect 18732 20468 18788 20478
rect 18508 20130 18564 20142
rect 18508 20078 18510 20130
rect 18562 20078 18564 20130
rect 18172 18286 18174 18338
rect 18226 18286 18228 18338
rect 18172 18228 18228 18286
rect 18172 18162 18228 18172
rect 18284 20018 18340 20030
rect 18284 19966 18286 20018
rect 18338 19966 18340 20018
rect 18284 17780 18340 19966
rect 18508 19908 18564 20078
rect 18620 20132 18676 20142
rect 18620 20038 18676 20076
rect 18508 19842 18564 19852
rect 18508 18452 18564 18462
rect 18564 18396 18676 18452
rect 18508 18358 18564 18396
rect 18284 17714 18340 17724
rect 18620 17668 18676 18396
rect 18620 17574 18676 17612
rect 18508 17444 18564 17454
rect 18732 17444 18788 20412
rect 18844 20244 18900 20750
rect 18956 20580 19012 23772
rect 19180 23380 19236 23390
rect 19628 23380 19684 24108
rect 19740 24098 19796 24108
rect 20412 24164 20468 26238
rect 20636 26292 20692 26302
rect 21084 26292 21140 26302
rect 21196 26292 21252 26798
rect 21308 26516 21364 27804
rect 21420 27746 21476 31892
rect 21756 28642 21812 28654
rect 21756 28590 21758 28642
rect 21810 28590 21812 28642
rect 21756 27860 21812 28590
rect 24668 28532 24724 28542
rect 21756 27766 21812 27804
rect 22316 27860 22372 27870
rect 21420 27694 21422 27746
rect 21474 27694 21476 27746
rect 21420 26962 21476 27694
rect 22316 27074 22372 27804
rect 22540 27748 22596 27758
rect 24668 27748 24724 28476
rect 22540 27654 22596 27692
rect 24444 27746 24724 27748
rect 24444 27694 24670 27746
rect 24722 27694 24724 27746
rect 24444 27692 24724 27694
rect 22316 27022 22318 27074
rect 22370 27022 22372 27074
rect 21420 26910 21422 26962
rect 21474 26910 21476 26962
rect 21420 26898 21476 26910
rect 21532 26964 21588 26974
rect 21532 26870 21588 26908
rect 22316 26852 22372 27022
rect 22988 26964 23044 26974
rect 22316 26786 22372 26796
rect 22652 26962 23044 26964
rect 22652 26910 22990 26962
rect 23042 26910 23044 26962
rect 22652 26908 23044 26910
rect 21420 26516 21476 26526
rect 21308 26514 21476 26516
rect 21308 26462 21422 26514
rect 21474 26462 21476 26514
rect 21308 26460 21476 26462
rect 21420 26450 21476 26460
rect 22652 26514 22708 26908
rect 22988 26898 23044 26908
rect 23548 26964 23604 26974
rect 23324 26516 23380 26526
rect 22652 26462 22654 26514
rect 22706 26462 22708 26514
rect 22652 26450 22708 26462
rect 22764 26514 23380 26516
rect 22764 26462 23326 26514
rect 23378 26462 23380 26514
rect 22764 26460 23380 26462
rect 20692 26236 21028 26292
rect 20636 26198 20692 26236
rect 20412 24098 20468 24108
rect 20748 24722 20804 24734
rect 20748 24670 20750 24722
rect 20802 24670 20804 24722
rect 20748 23828 20804 24670
rect 20748 23762 20804 23772
rect 20972 24498 21028 26236
rect 21084 26290 21252 26292
rect 21084 26238 21086 26290
rect 21138 26238 21252 26290
rect 21084 26236 21252 26238
rect 21308 26292 21364 26302
rect 21084 26226 21140 26236
rect 21196 24836 21252 24846
rect 21196 24722 21252 24780
rect 21308 24834 21364 26236
rect 22540 26292 22596 26302
rect 22764 26292 22820 26460
rect 23324 26450 23380 26460
rect 23436 26516 23492 26526
rect 23436 26422 23492 26460
rect 23548 26514 23604 26908
rect 23548 26462 23550 26514
rect 23602 26462 23604 26514
rect 23548 26450 23604 26462
rect 24332 26964 24388 26974
rect 24332 26514 24388 26908
rect 24332 26462 24334 26514
rect 24386 26462 24388 26514
rect 24332 26450 24388 26462
rect 24444 26514 24500 27692
rect 24668 27682 24724 27692
rect 25116 27186 25172 37996
rect 26236 37940 26292 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 26236 37874 26292 37884
rect 27468 37940 27524 37950
rect 27468 37846 27524 37884
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 25228 37266 25284 37278
rect 25228 37214 25230 37266
rect 25282 37214 25284 37266
rect 25228 28532 25284 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 25228 28466 25284 28476
rect 25116 27134 25118 27186
rect 25170 27134 25172 27186
rect 24444 26462 24446 26514
rect 24498 26462 24500 26514
rect 24444 26450 24500 26462
rect 24556 27076 24612 27086
rect 24556 26514 24612 27020
rect 24556 26462 24558 26514
rect 24610 26462 24612 26514
rect 24556 26450 24612 26462
rect 25116 26516 25172 27134
rect 25116 26450 25172 26460
rect 25340 27746 25396 27758
rect 25340 27694 25342 27746
rect 25394 27694 25396 27746
rect 25340 26852 25396 27694
rect 25452 27748 25508 27758
rect 25452 27298 25508 27692
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25452 27246 25454 27298
rect 25506 27246 25508 27298
rect 25452 27234 25508 27246
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 37660 27074 37716 27086
rect 37660 27022 37662 27074
rect 37714 27022 37716 27074
rect 25564 26964 25620 26974
rect 25564 26870 25620 26908
rect 22540 26290 22820 26292
rect 22540 26238 22542 26290
rect 22594 26238 22820 26290
rect 22540 26236 22820 26238
rect 23100 26290 23156 26302
rect 23100 26238 23102 26290
rect 23154 26238 23156 26290
rect 22540 26226 22596 26236
rect 23100 25956 23156 26238
rect 23212 26292 23268 26302
rect 23212 26198 23268 26236
rect 24108 26290 24164 26302
rect 24108 26238 24110 26290
rect 24162 26238 24164 26290
rect 23100 25900 23268 25956
rect 23212 25284 23268 25900
rect 21308 24782 21310 24834
rect 21362 24782 21364 24834
rect 21308 24770 21364 24782
rect 21420 24948 21476 24958
rect 21196 24670 21198 24722
rect 21250 24670 21252 24722
rect 21196 24658 21252 24670
rect 20972 24446 20974 24498
rect 21026 24446 21028 24498
rect 20076 23716 20132 23726
rect 20132 23660 20244 23716
rect 20076 23650 20132 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23380 20244 23660
rect 19180 23378 19684 23380
rect 19180 23326 19182 23378
rect 19234 23326 19684 23378
rect 19180 23324 19684 23326
rect 19180 23314 19236 23324
rect 19068 23266 19124 23278
rect 19068 23214 19070 23266
rect 19122 23214 19124 23266
rect 19068 22372 19124 23214
rect 19628 23266 19684 23324
rect 19628 23214 19630 23266
rect 19682 23214 19684 23266
rect 19628 23202 19684 23214
rect 20076 23324 20244 23380
rect 19516 23154 19572 23166
rect 19516 23102 19518 23154
rect 19570 23102 19572 23154
rect 19068 22316 19348 22372
rect 19180 22146 19236 22158
rect 19180 22094 19182 22146
rect 19234 22094 19236 22146
rect 19180 20804 19236 22094
rect 19180 20738 19236 20748
rect 19180 20580 19236 20590
rect 18956 20578 19236 20580
rect 18956 20526 19182 20578
rect 19234 20526 19236 20578
rect 18956 20524 19236 20526
rect 18844 20178 18900 20188
rect 19068 20242 19124 20524
rect 19180 20514 19236 20524
rect 19292 20468 19348 22316
rect 19292 20402 19348 20412
rect 19516 20468 19572 23102
rect 19852 23156 19908 23166
rect 19852 23062 19908 23100
rect 20076 23154 20132 23324
rect 20076 23102 20078 23154
rect 20130 23102 20132 23154
rect 20076 23090 20132 23102
rect 20412 23154 20468 23166
rect 20412 23102 20414 23154
rect 20466 23102 20468 23154
rect 20412 23044 20468 23102
rect 20412 22978 20468 22988
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19852 21812 19908 21822
rect 19628 21364 19684 21374
rect 19628 20802 19684 21308
rect 19628 20750 19630 20802
rect 19682 20750 19684 20802
rect 19628 20738 19684 20750
rect 19852 21028 19908 21756
rect 19852 20802 19908 20972
rect 20300 21476 20356 21486
rect 19852 20750 19854 20802
rect 19906 20750 19908 20802
rect 19852 20738 19908 20750
rect 20188 20804 20244 20814
rect 20188 20710 20244 20748
rect 20076 20692 20132 20702
rect 19964 20580 20020 20618
rect 20076 20598 20132 20636
rect 19964 20514 20020 20524
rect 19516 20402 19572 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20300 20356 20356 21420
rect 19836 20346 20100 20356
rect 20188 20300 20356 20356
rect 20636 21028 20692 21038
rect 19068 20190 19070 20242
rect 19122 20190 19124 20242
rect 19068 20178 19124 20190
rect 19964 20244 20020 20254
rect 19964 20150 20020 20188
rect 19404 20132 19460 20142
rect 19292 20018 19348 20030
rect 19292 19966 19294 20018
rect 19346 19966 19348 20018
rect 19292 19348 19348 19966
rect 19404 19796 19460 20076
rect 19404 19730 19460 19740
rect 19516 20018 19572 20030
rect 19516 19966 19518 20018
rect 19570 19966 19572 20018
rect 19292 19282 19348 19292
rect 19516 19124 19572 19966
rect 18844 19068 19572 19124
rect 19628 20020 19684 20030
rect 18844 18562 18900 19068
rect 18844 18510 18846 18562
rect 18898 18510 18900 18562
rect 18844 18340 18900 18510
rect 18844 18274 18900 18284
rect 19180 17890 19236 19068
rect 19628 18676 19684 19964
rect 19740 20018 19796 20030
rect 19740 19966 19742 20018
rect 19794 19966 19796 20018
rect 19740 19012 19796 19966
rect 20076 20020 20132 20030
rect 20076 19926 20132 19964
rect 20188 19796 20244 20300
rect 20524 20132 20580 20142
rect 20412 20130 20580 20132
rect 20412 20078 20526 20130
rect 20578 20078 20580 20130
rect 20412 20076 20580 20078
rect 20412 19908 20468 20076
rect 20524 20066 20580 20076
rect 20636 20130 20692 20972
rect 20972 20804 21028 24446
rect 21084 23156 21140 23166
rect 21084 23062 21140 23100
rect 20972 20738 21028 20748
rect 21420 20244 21476 24892
rect 22540 24948 22596 24958
rect 22540 24854 22596 24892
rect 22316 24836 22372 24846
rect 22316 24742 22372 24780
rect 22204 24722 22260 24734
rect 22204 24670 22206 24722
rect 22258 24670 22260 24722
rect 22204 24612 22260 24670
rect 22204 24546 22260 24556
rect 22540 23826 22596 23838
rect 22540 23774 22542 23826
rect 22594 23774 22596 23826
rect 22204 23716 22260 23726
rect 22204 23622 22260 23660
rect 22428 23714 22484 23726
rect 22428 23662 22430 23714
rect 22482 23662 22484 23714
rect 22428 23268 22484 23662
rect 22428 23202 22484 23212
rect 21980 22370 22036 22382
rect 21980 22318 21982 22370
rect 22034 22318 22036 22370
rect 21868 21812 21924 21822
rect 21532 21588 21588 21598
rect 21532 20802 21588 21532
rect 21532 20750 21534 20802
rect 21586 20750 21588 20802
rect 21532 20468 21588 20750
rect 21532 20402 21588 20412
rect 21644 21028 21700 21038
rect 20636 20078 20638 20130
rect 20690 20078 20692 20130
rect 20636 20066 20692 20078
rect 21308 20188 21476 20244
rect 20412 19842 20468 19852
rect 20076 19740 20244 19796
rect 20524 19794 20580 19806
rect 20524 19742 20526 19794
rect 20578 19742 20580 19794
rect 20076 19234 20132 19740
rect 20076 19182 20078 19234
rect 20130 19182 20132 19234
rect 20076 19170 20132 19182
rect 20188 19348 20244 19358
rect 19740 18946 19796 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19964 18676 20020 18686
rect 20188 18676 20244 19292
rect 19628 18674 19908 18676
rect 19628 18622 19630 18674
rect 19682 18622 19908 18674
rect 19628 18620 19908 18622
rect 19628 18610 19684 18620
rect 19180 17838 19182 17890
rect 19234 17838 19236 17890
rect 19180 17826 19236 17838
rect 18508 17442 18788 17444
rect 18508 17390 18510 17442
rect 18562 17390 18788 17442
rect 18508 17388 18788 17390
rect 18508 17378 18564 17388
rect 18060 16230 18116 16268
rect 17724 16098 17892 16100
rect 17724 16046 17726 16098
rect 17778 16046 17892 16098
rect 17724 16044 17892 16046
rect 17724 16034 17780 16044
rect 18396 15988 18452 15998
rect 17612 15876 17668 15886
rect 18172 15876 18228 15886
rect 17276 15810 17332 15820
rect 17500 15874 17668 15876
rect 17500 15822 17614 15874
rect 17666 15822 17668 15874
rect 17500 15820 17668 15822
rect 17388 15428 17444 15438
rect 16380 15262 16382 15314
rect 16434 15262 16436 15314
rect 16380 15250 16436 15262
rect 16604 15316 16660 15326
rect 16604 15222 16660 15260
rect 16716 15204 16772 15242
rect 16716 15138 16772 15148
rect 16268 15092 16324 15102
rect 15372 15090 16324 15092
rect 15372 15038 16270 15090
rect 16322 15038 16324 15090
rect 15372 15036 16324 15038
rect 15372 14642 15428 15036
rect 16268 15026 16324 15036
rect 15372 14590 15374 14642
rect 15426 14590 15428 14642
rect 15372 14578 15428 14590
rect 17388 14644 17444 15372
rect 17500 15316 17556 15820
rect 17612 15810 17668 15820
rect 17724 15874 18228 15876
rect 17724 15822 18174 15874
rect 18226 15822 18228 15874
rect 17724 15820 18228 15822
rect 17500 15092 17556 15260
rect 17612 15316 17668 15326
rect 17724 15316 17780 15820
rect 18172 15810 18228 15820
rect 18284 15874 18340 15886
rect 18284 15822 18286 15874
rect 18338 15822 18340 15874
rect 18284 15764 18340 15822
rect 18284 15698 18340 15708
rect 18396 15540 18452 15932
rect 18732 15876 18788 17388
rect 18732 15810 18788 15820
rect 18956 17780 19012 17790
rect 17948 15484 18452 15540
rect 17948 15426 18004 15484
rect 17948 15374 17950 15426
rect 18002 15374 18004 15426
rect 17948 15362 18004 15374
rect 18732 15428 18788 15438
rect 17612 15314 17780 15316
rect 17612 15262 17614 15314
rect 17666 15262 17780 15314
rect 17612 15260 17780 15262
rect 18172 15316 18228 15326
rect 18508 15316 18564 15326
rect 18172 15314 18340 15316
rect 18172 15262 18174 15314
rect 18226 15262 18340 15314
rect 18172 15260 18340 15262
rect 17612 15250 17668 15260
rect 18172 15250 18228 15260
rect 18060 15202 18116 15214
rect 18060 15150 18062 15202
rect 18114 15150 18116 15202
rect 17612 15092 17668 15102
rect 17500 15090 17668 15092
rect 17500 15038 17614 15090
rect 17666 15038 17668 15090
rect 17500 15036 17668 15038
rect 17612 15026 17668 15036
rect 17500 14644 17556 14654
rect 17388 14642 17556 14644
rect 17388 14590 17502 14642
rect 17554 14590 17556 14642
rect 17388 14588 17556 14590
rect 14700 14438 14756 14476
rect 16380 14532 16436 14542
rect 16380 13972 16436 14476
rect 16828 13972 16884 13982
rect 16380 13970 16828 13972
rect 16380 13918 16382 13970
rect 16434 13918 16828 13970
rect 16380 13916 16828 13918
rect 16380 13906 16436 13916
rect 16828 13878 16884 13916
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 17388 8428 17444 14588
rect 17500 14578 17556 14588
rect 17948 14532 18004 14542
rect 17948 14438 18004 14476
rect 17500 13972 17556 13982
rect 17500 13746 17556 13916
rect 18060 13860 18116 15150
rect 18284 15148 18340 15260
rect 18508 15148 18564 15260
rect 18732 15314 18788 15372
rect 18732 15262 18734 15314
rect 18786 15262 18788 15314
rect 18732 15250 18788 15262
rect 18284 15092 18564 15148
rect 18620 15204 18676 15242
rect 18956 15148 19012 17724
rect 19852 17666 19908 18620
rect 19964 18674 20188 18676
rect 19964 18622 19966 18674
rect 20018 18622 20188 18674
rect 19964 18620 20188 18622
rect 19964 18610 20020 18620
rect 20188 18582 20244 18620
rect 20412 19236 20468 19246
rect 20300 18452 20356 18462
rect 20300 18358 20356 18396
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17602 19908 17614
rect 20188 17556 20244 17566
rect 20412 17556 20468 19180
rect 20188 17554 20468 17556
rect 20188 17502 20190 17554
rect 20242 17502 20468 17554
rect 20188 17500 20468 17502
rect 20188 17490 20244 17500
rect 19516 17444 19572 17454
rect 19516 17350 19572 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20076 17108 20132 17118
rect 19292 16884 19348 16894
rect 19180 15988 19236 15998
rect 18620 15138 18676 15148
rect 18844 15092 19012 15148
rect 19068 15932 19180 15988
rect 18284 14418 18340 15092
rect 18732 14756 18788 14766
rect 18844 14756 18900 15092
rect 18732 14754 18900 14756
rect 18732 14702 18734 14754
rect 18786 14702 18900 14754
rect 18732 14700 18900 14702
rect 18956 14756 19012 14766
rect 19068 14756 19124 15932
rect 19180 15894 19236 15932
rect 19180 15316 19236 15326
rect 19292 15316 19348 16828
rect 19404 16100 19460 16110
rect 19404 16006 19460 16044
rect 19180 15314 19348 15316
rect 19180 15262 19182 15314
rect 19234 15262 19348 15314
rect 19180 15260 19348 15262
rect 19404 15876 19460 15886
rect 20076 15876 20132 17052
rect 20524 17108 20580 19742
rect 21308 19460 21364 20188
rect 21532 20130 21588 20142
rect 21532 20078 21534 20130
rect 21586 20078 21588 20130
rect 20748 19404 21364 19460
rect 21420 20020 21476 20030
rect 21420 19460 21476 19964
rect 21532 19796 21588 20078
rect 21532 19730 21588 19740
rect 21420 19404 21588 19460
rect 20636 18562 20692 18574
rect 20636 18510 20638 18562
rect 20690 18510 20692 18562
rect 20636 18340 20692 18510
rect 20636 18274 20692 18284
rect 20748 17556 20804 19404
rect 21196 19234 21252 19246
rect 21196 19182 21198 19234
rect 21250 19182 21252 19234
rect 20972 18676 21028 18686
rect 20972 18562 21028 18620
rect 20972 18510 20974 18562
rect 21026 18510 21028 18562
rect 20972 18452 21028 18510
rect 21084 18564 21140 18574
rect 21196 18564 21252 19182
rect 21308 19236 21364 19404
rect 21420 19236 21476 19246
rect 21308 19234 21476 19236
rect 21308 19182 21422 19234
rect 21474 19182 21476 19234
rect 21308 19180 21476 19182
rect 21420 19170 21476 19180
rect 21308 18676 21364 18686
rect 21532 18676 21588 19404
rect 21308 18674 21588 18676
rect 21308 18622 21310 18674
rect 21362 18622 21588 18674
rect 21308 18620 21588 18622
rect 21644 19234 21700 20972
rect 21868 20690 21924 21756
rect 21980 21476 22036 22318
rect 22540 21812 22596 23774
rect 23212 23826 23268 25228
rect 24108 25284 24164 26238
rect 24108 25218 24164 25228
rect 24220 26290 24276 26302
rect 24220 26238 24222 26290
rect 24274 26238 24276 26290
rect 23212 23774 23214 23826
rect 23266 23774 23268 23826
rect 23212 23762 23268 23774
rect 23772 24948 23828 24958
rect 22540 21746 22596 21756
rect 22876 23714 22932 23726
rect 22876 23662 22878 23714
rect 22930 23662 22932 23714
rect 21980 21410 22036 21420
rect 22876 21028 22932 23662
rect 23548 23380 23604 23390
rect 23212 23268 23268 23278
rect 23212 23042 23268 23212
rect 23548 23266 23604 23324
rect 23548 23214 23550 23266
rect 23602 23214 23604 23266
rect 23548 23202 23604 23214
rect 23772 23378 23828 24892
rect 24220 24612 24276 26238
rect 25340 26292 25396 26796
rect 26012 26852 26068 26862
rect 26012 26758 26068 26796
rect 25452 26292 25508 26302
rect 25340 26290 25508 26292
rect 25340 26238 25454 26290
rect 25506 26238 25508 26290
rect 25340 26236 25508 26238
rect 25116 25284 25172 25294
rect 25452 25284 25508 26236
rect 26236 26180 26292 26190
rect 26012 26178 26292 26180
rect 26012 26126 26238 26178
rect 26290 26126 26292 26178
rect 26012 26124 26292 26126
rect 26012 25618 26068 26124
rect 26236 26114 26292 26124
rect 27244 26180 27300 26190
rect 26012 25566 26014 25618
rect 26066 25566 26068 25618
rect 26012 25554 26068 25566
rect 26572 25508 26628 25518
rect 27020 25508 27076 25518
rect 26572 25506 27076 25508
rect 26572 25454 26574 25506
rect 26626 25454 27022 25506
rect 27074 25454 27076 25506
rect 26572 25452 27076 25454
rect 26572 25442 26628 25452
rect 27020 25442 27076 25452
rect 27244 25394 27300 26124
rect 28364 26180 28420 26190
rect 28364 26086 28420 26124
rect 37660 26180 37716 27022
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 37660 26114 37716 26124
rect 27356 26068 27412 26078
rect 27356 25508 27412 26012
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 27804 25508 27860 25518
rect 27356 25506 27860 25508
rect 27356 25454 27358 25506
rect 27410 25454 27806 25506
rect 27858 25454 27860 25506
rect 27356 25452 27860 25454
rect 27356 25442 27412 25452
rect 27244 25342 27246 25394
rect 27298 25342 27300 25394
rect 27244 25330 27300 25342
rect 25116 25282 25508 25284
rect 25116 25230 25118 25282
rect 25170 25230 25508 25282
rect 25116 25228 25508 25230
rect 25900 25282 25956 25294
rect 25900 25230 25902 25282
rect 25954 25230 25956 25282
rect 25116 25218 25172 25228
rect 24220 24546 24276 24556
rect 25228 23716 25284 25228
rect 25900 24948 25956 25230
rect 26124 25284 26180 25294
rect 26124 24948 26180 25228
rect 26124 24892 26628 24948
rect 25900 24882 25956 24892
rect 25676 23938 25732 23950
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25340 23716 25396 23726
rect 25676 23716 25732 23886
rect 25228 23714 25732 23716
rect 25228 23662 25342 23714
rect 25394 23662 25732 23714
rect 25228 23660 25732 23662
rect 26460 23826 26516 23838
rect 26460 23774 26462 23826
rect 26514 23774 26516 23826
rect 23772 23326 23774 23378
rect 23826 23326 23828 23378
rect 23212 22990 23214 23042
rect 23266 22990 23268 23042
rect 23212 22978 23268 22990
rect 22876 20962 22932 20972
rect 23660 22930 23716 22942
rect 23660 22878 23662 22930
rect 23714 22878 23716 22930
rect 22204 20916 22260 20926
rect 22204 20802 22260 20860
rect 23660 20914 23716 22878
rect 23660 20862 23662 20914
rect 23714 20862 23716 20914
rect 23660 20850 23716 20862
rect 22204 20750 22206 20802
rect 22258 20750 22260 20802
rect 22204 20738 22260 20750
rect 22876 20802 22932 20814
rect 22876 20750 22878 20802
rect 22930 20750 22932 20802
rect 21868 20638 21870 20690
rect 21922 20638 21924 20690
rect 21868 20626 21924 20638
rect 22316 20692 22372 20702
rect 21868 20468 21924 20478
rect 21756 20356 21812 20366
rect 21756 20130 21812 20300
rect 21756 20078 21758 20130
rect 21810 20078 21812 20130
rect 21756 20066 21812 20078
rect 21644 19182 21646 19234
rect 21698 19182 21700 19234
rect 21308 18610 21364 18620
rect 21140 18508 21252 18564
rect 21084 18470 21140 18508
rect 20972 18386 21028 18396
rect 21644 18340 21700 19182
rect 21868 19236 21924 20412
rect 21980 20132 22036 20142
rect 21980 20038 22036 20076
rect 22092 20130 22148 20142
rect 22092 20078 22094 20130
rect 22146 20078 22148 20130
rect 22092 20020 22148 20078
rect 22316 20130 22372 20636
rect 22316 20078 22318 20130
rect 22370 20078 22372 20130
rect 22316 20066 22372 20078
rect 22540 20580 22596 20590
rect 22092 19954 22148 19964
rect 22204 19236 22260 19246
rect 22540 19236 22596 20524
rect 22876 20244 22932 20750
rect 22876 20178 22932 20188
rect 23660 20244 23716 20254
rect 21924 19234 22260 19236
rect 21924 19182 22206 19234
rect 22258 19182 22260 19234
rect 21924 19180 22260 19182
rect 21868 19142 21924 19180
rect 22204 19170 22260 19180
rect 22316 19180 22596 19236
rect 22316 19012 22372 19180
rect 22540 19012 22596 19022
rect 21644 18274 21700 18284
rect 22204 18956 22372 19012
rect 22428 18956 22540 19012
rect 20524 17042 20580 17052
rect 20636 17500 20804 17556
rect 22204 17556 22260 18956
rect 20076 15820 20244 15876
rect 19180 15250 19236 15260
rect 19404 15148 19460 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19964 15540 20020 15550
rect 20188 15540 20244 15820
rect 18956 14754 19124 14756
rect 18956 14702 18958 14754
rect 19010 14702 19124 14754
rect 18956 14700 19124 14702
rect 19180 15092 19460 15148
rect 19516 15316 19572 15326
rect 18732 14690 18788 14700
rect 18956 14690 19012 14700
rect 19180 14642 19236 15092
rect 19404 14644 19460 14654
rect 19180 14590 19182 14642
rect 19234 14590 19236 14642
rect 19180 14578 19236 14590
rect 19292 14642 19460 14644
rect 19292 14590 19406 14642
rect 19458 14590 19460 14642
rect 19292 14588 19460 14590
rect 18284 14366 18286 14418
rect 18338 14366 18340 14418
rect 18284 14354 18340 14366
rect 18172 13860 18228 13870
rect 18060 13858 18228 13860
rect 18060 13806 18174 13858
rect 18226 13806 18228 13858
rect 18060 13804 18228 13806
rect 18172 13794 18228 13804
rect 17500 13694 17502 13746
rect 17554 13694 17556 13746
rect 17500 13076 17556 13694
rect 19292 13524 19348 14588
rect 19404 14578 19460 14588
rect 19404 14420 19460 14430
rect 19516 14420 19572 15260
rect 19404 14418 19572 14420
rect 19404 14366 19406 14418
rect 19458 14366 19572 14418
rect 19404 14364 19572 14366
rect 19404 14354 19460 14364
rect 19628 14308 19684 14318
rect 19964 14308 20020 15484
rect 20076 15484 20244 15540
rect 20076 15426 20132 15484
rect 20076 15374 20078 15426
rect 20130 15374 20132 15426
rect 20076 15362 20132 15374
rect 20300 15316 20356 15326
rect 20300 15222 20356 15260
rect 20524 15316 20580 15326
rect 20636 15316 20692 17500
rect 21532 17444 21588 17454
rect 20524 15314 20692 15316
rect 20524 15262 20526 15314
rect 20578 15262 20692 15314
rect 20524 15260 20692 15262
rect 20748 17332 20804 17342
rect 20748 15314 20804 17276
rect 21196 17108 21252 17118
rect 21196 17014 21252 17052
rect 21420 17108 21476 17118
rect 21420 15988 21476 17052
rect 21532 16994 21588 17388
rect 21532 16942 21534 16994
rect 21586 16942 21588 16994
rect 21532 16930 21588 16942
rect 21644 16994 21700 17006
rect 21644 16942 21646 16994
rect 21698 16942 21700 16994
rect 21644 16772 21700 16942
rect 22204 16884 22260 17500
rect 22316 17666 22372 17678
rect 22316 17614 22318 17666
rect 22370 17614 22372 17666
rect 22316 17444 22372 17614
rect 22316 17378 22372 17388
rect 22428 17332 22484 18956
rect 22540 18918 22596 18956
rect 23660 19010 23716 20188
rect 23772 19908 23828 23326
rect 23996 23266 24052 23278
rect 23996 23214 23998 23266
rect 24050 23214 24052 23266
rect 23884 21586 23940 21598
rect 23884 21534 23886 21586
rect 23938 21534 23940 21586
rect 23884 20580 23940 21534
rect 23996 21474 24052 23214
rect 24444 23044 24500 23054
rect 24444 22260 24500 22988
rect 24444 22194 24500 22204
rect 25340 22260 25396 23660
rect 26348 23380 26404 23390
rect 26460 23380 26516 23774
rect 26348 23378 26516 23380
rect 26348 23326 26350 23378
rect 26402 23326 26516 23378
rect 26348 23324 26516 23326
rect 26348 23314 26404 23324
rect 26236 23156 26292 23166
rect 26460 23156 26516 23166
rect 26572 23156 26628 24892
rect 27356 24052 27412 24062
rect 27356 23378 27412 23996
rect 27356 23326 27358 23378
rect 27410 23326 27412 23378
rect 27356 23314 27412 23326
rect 27468 23380 27524 25452
rect 27804 25442 27860 25452
rect 37660 24722 37716 24734
rect 37660 24670 37662 24722
rect 37714 24670 37716 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 28588 24052 28644 24062
rect 28588 23958 28644 23996
rect 37660 24052 37716 24670
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 40012 24276 40068 24446
rect 40012 24210 40068 24220
rect 37660 23986 37716 23996
rect 27916 23380 27972 23390
rect 27468 23378 27972 23380
rect 27468 23326 27918 23378
rect 27970 23326 27972 23378
rect 27468 23324 27972 23326
rect 27468 23266 27524 23324
rect 27916 23314 27972 23324
rect 27468 23214 27470 23266
rect 27522 23214 27524 23266
rect 27468 23202 27524 23214
rect 26236 23154 26404 23156
rect 26236 23102 26238 23154
rect 26290 23102 26404 23154
rect 26236 23100 26404 23102
rect 26236 23090 26292 23100
rect 26348 22484 26404 23100
rect 26460 23154 26628 23156
rect 26460 23102 26462 23154
rect 26514 23102 26628 23154
rect 26460 23100 26628 23102
rect 26908 23156 26964 23166
rect 27132 23156 27188 23166
rect 26908 23154 27188 23156
rect 26908 23102 26910 23154
rect 26962 23102 27134 23154
rect 27186 23102 27188 23154
rect 26908 23100 27188 23102
rect 26460 23090 26516 23100
rect 26908 23090 26964 23100
rect 27132 23090 27188 23100
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 26348 22428 26852 22484
rect 25340 22194 25396 22204
rect 25788 22260 25844 22270
rect 23996 21422 23998 21474
rect 24050 21422 24052 21474
rect 23996 21410 24052 21422
rect 24108 21812 24164 21822
rect 23884 20514 23940 20524
rect 24108 20244 24164 21756
rect 24332 21698 24388 21710
rect 24332 21646 24334 21698
rect 24386 21646 24388 21698
rect 24332 21252 24388 21646
rect 25788 21586 25844 22204
rect 25788 21534 25790 21586
rect 25842 21534 25844 21586
rect 24332 21186 24388 21196
rect 25452 21476 25508 21486
rect 25788 21476 25844 21534
rect 25452 21474 25844 21476
rect 25452 21422 25454 21474
rect 25506 21422 25844 21474
rect 25452 21420 25844 21422
rect 24108 20178 24164 20188
rect 24332 20916 24388 20926
rect 24332 20130 24388 20860
rect 25228 20916 25284 20926
rect 25452 20916 25508 21420
rect 25284 20860 25508 20916
rect 25788 21252 25844 21262
rect 25788 20914 25844 21196
rect 25788 20862 25790 20914
rect 25842 20862 25844 20914
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24332 20066 24388 20078
rect 24668 20132 24724 20142
rect 24668 20038 24724 20076
rect 23772 19852 24388 19908
rect 24332 19122 24388 19852
rect 24332 19070 24334 19122
rect 24386 19070 24388 19122
rect 24332 19058 24388 19070
rect 24556 19796 24612 19806
rect 24556 19122 24612 19740
rect 24556 19070 24558 19122
rect 24610 19070 24612 19122
rect 24556 19058 24612 19070
rect 24780 19346 24836 19358
rect 24780 19294 24782 19346
rect 24834 19294 24836 19346
rect 24780 19124 24836 19294
rect 25228 19236 25284 20860
rect 25788 20850 25844 20862
rect 25900 20748 26180 20804
rect 25900 20242 25956 20748
rect 26124 20692 26180 20748
rect 26236 20692 26292 20702
rect 26124 20690 26292 20692
rect 26124 20638 26238 20690
rect 26290 20638 26292 20690
rect 26124 20636 26292 20638
rect 26236 20626 26292 20636
rect 26348 20692 26404 20702
rect 26348 20598 26404 20636
rect 25900 20190 25902 20242
rect 25954 20190 25956 20242
rect 25900 20178 25956 20190
rect 26012 20578 26068 20590
rect 26012 20526 26014 20578
rect 26066 20526 26068 20578
rect 25340 20132 25396 20142
rect 25340 20038 25396 20076
rect 25788 20130 25844 20142
rect 25788 20078 25790 20130
rect 25842 20078 25844 20130
rect 25564 20018 25620 20030
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 25228 19234 25396 19236
rect 25228 19182 25230 19234
rect 25282 19182 25396 19234
rect 25228 19180 25396 19182
rect 25228 19170 25284 19180
rect 24780 19058 24836 19068
rect 23660 18958 23662 19010
rect 23714 18958 23716 19010
rect 22652 18452 22708 18462
rect 22428 17266 22484 17276
rect 22540 18340 22596 18350
rect 22540 17220 22596 18284
rect 22540 17106 22596 17164
rect 22540 17054 22542 17106
rect 22594 17054 22596 17106
rect 22540 17042 22596 17054
rect 22652 16996 22708 18396
rect 23660 18452 23716 18958
rect 23660 18386 23716 18396
rect 23996 19010 24052 19022
rect 23996 18958 23998 19010
rect 24050 18958 24052 19010
rect 23996 17892 24052 18958
rect 24220 19012 24276 19022
rect 24220 18918 24276 18956
rect 23996 17826 24052 17836
rect 24668 18452 24724 18462
rect 24668 18338 24724 18396
rect 25340 18452 25396 19180
rect 25564 19012 25620 19966
rect 25788 19348 25844 20078
rect 25788 19282 25844 19292
rect 25900 19124 25956 19134
rect 25900 19030 25956 19068
rect 25564 18946 25620 18956
rect 25340 18358 25396 18396
rect 26012 18450 26068 20526
rect 26460 20468 26516 22428
rect 26796 22370 26852 22428
rect 26796 22318 26798 22370
rect 26850 22318 26852 22370
rect 26796 22306 26852 22318
rect 27020 22482 27076 22494
rect 27020 22430 27022 22482
rect 27074 22430 27076 22482
rect 27020 21924 27076 22430
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 37884 22370 37940 22382
rect 37884 22318 37886 22370
rect 37938 22318 37940 22370
rect 26908 21868 27076 21924
rect 27132 22146 27188 22158
rect 27132 22094 27134 22146
rect 27186 22094 27188 22146
rect 26572 21476 26628 21486
rect 26572 21474 26852 21476
rect 26572 21422 26574 21474
rect 26626 21422 26852 21474
rect 26572 21420 26852 21422
rect 26572 21410 26628 21420
rect 26796 21026 26852 21420
rect 26796 20974 26798 21026
rect 26850 20974 26852 21026
rect 26796 20962 26852 20974
rect 26908 20804 26964 21868
rect 26796 20748 26964 20804
rect 26124 20412 26516 20468
rect 26684 20690 26740 20702
rect 26684 20638 26686 20690
rect 26738 20638 26740 20690
rect 26124 20132 26180 20412
rect 26684 20356 26740 20638
rect 26796 20690 26852 20748
rect 26796 20638 26798 20690
rect 26850 20638 26852 20690
rect 26796 20626 26852 20638
rect 26684 20290 26740 20300
rect 26124 20038 26180 20076
rect 26348 20244 26404 20254
rect 26348 20130 26404 20188
rect 27132 20244 27188 22094
rect 27356 22146 27412 22158
rect 27356 22094 27358 22146
rect 27410 22094 27412 22146
rect 27356 21476 27412 22094
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 27356 21410 27412 21420
rect 28700 21476 28756 21486
rect 28700 21382 28756 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 37884 21028 37940 22318
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 40012 21588 40068 21598
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 37884 20962 37940 20972
rect 27356 20916 27412 20926
rect 27356 20822 27412 20860
rect 27132 20178 27188 20188
rect 26348 20078 26350 20130
rect 26402 20078 26404 20130
rect 26348 20066 26404 20078
rect 26572 20130 26628 20142
rect 26572 20078 26574 20130
rect 26626 20078 26628 20130
rect 26236 19796 26292 19806
rect 26236 19702 26292 19740
rect 26572 19348 26628 20078
rect 37660 20018 37716 20030
rect 37660 19966 37662 20018
rect 37714 19966 37716 20018
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 37660 19460 37716 19966
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 37660 19394 37716 19404
rect 26572 19282 26628 19292
rect 28028 19348 28084 19358
rect 28028 19254 28084 19292
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 37660 19236 37716 19246
rect 37660 19142 37716 19180
rect 26012 18398 26014 18450
rect 26066 18398 26068 18450
rect 26012 18386 26068 18398
rect 28140 19124 28196 19134
rect 24668 18286 24670 18338
rect 24722 18286 24724 18338
rect 22652 16902 22708 16940
rect 22764 17554 22820 17566
rect 22764 17502 22766 17554
rect 22818 17502 22820 17554
rect 22316 16884 22372 16894
rect 22204 16828 22316 16884
rect 22316 16790 22372 16828
rect 21644 16706 21700 16716
rect 21980 16770 22036 16782
rect 21980 16718 21982 16770
rect 22034 16718 22036 16770
rect 21420 15922 21476 15932
rect 21084 15540 21140 15550
rect 21084 15538 21812 15540
rect 21084 15486 21086 15538
rect 21138 15486 21812 15538
rect 21084 15484 21812 15486
rect 21084 15474 21140 15484
rect 20748 15262 20750 15314
rect 20802 15262 20804 15314
rect 20524 15250 20580 15260
rect 20748 15250 20804 15262
rect 20972 15314 21028 15326
rect 20972 15262 20974 15314
rect 21026 15262 21028 15314
rect 20972 14756 21028 15262
rect 20972 14690 21028 14700
rect 21308 15316 21364 15326
rect 20524 14418 20580 14430
rect 20524 14366 20526 14418
rect 20578 14366 20580 14418
rect 20412 14308 20468 14318
rect 19964 14252 20244 14308
rect 19628 14214 19684 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13636 20244 14252
rect 20412 14214 20468 14252
rect 20300 13636 20356 13646
rect 18620 13468 19348 13524
rect 19628 13634 20356 13636
rect 19628 13582 20302 13634
rect 20354 13582 20356 13634
rect 19628 13580 20356 13582
rect 17612 13076 17668 13086
rect 17500 13074 17892 13076
rect 17500 13022 17614 13074
rect 17666 13022 17892 13074
rect 17500 13020 17892 13022
rect 17612 13010 17668 13020
rect 17836 12962 17892 13020
rect 18620 13074 18676 13468
rect 18620 13022 18622 13074
rect 18674 13022 18676 13074
rect 18620 13010 18676 13022
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 17836 12898 17892 12910
rect 17388 8372 17780 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 17724 4338 17780 8372
rect 17724 4286 17726 4338
rect 17778 4286 17780 4338
rect 17724 4274 17780 4286
rect 17500 4116 17556 4126
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17500 800 17556 4060
rect 18732 4116 18788 4126
rect 18732 4022 18788 4060
rect 18172 3666 18228 3678
rect 18172 3614 18174 3666
rect 18226 3614 18228 3666
rect 18172 800 18228 3614
rect 19628 3556 19684 13580
rect 20300 13570 20356 13580
rect 20524 13076 20580 14366
rect 21084 13748 21140 13758
rect 21308 13748 21364 15260
rect 21756 13858 21812 15484
rect 21980 15428 22036 16718
rect 22428 16772 22484 16782
rect 22428 16678 22484 16716
rect 22764 16772 22820 17502
rect 23436 17556 23492 17566
rect 22876 17442 22932 17454
rect 22876 17390 22878 17442
rect 22930 17390 22932 17442
rect 22876 17108 22932 17390
rect 22988 17442 23044 17454
rect 22988 17390 22990 17442
rect 23042 17390 23044 17442
rect 22988 17108 23044 17390
rect 23100 17442 23156 17454
rect 23100 17390 23102 17442
rect 23154 17390 23156 17442
rect 23100 17332 23156 17390
rect 23100 17266 23156 17276
rect 22988 17052 23156 17108
rect 22876 17042 22932 17052
rect 22988 16884 23044 16894
rect 22988 16790 23044 16828
rect 22764 16706 22820 16716
rect 23100 16212 23156 17052
rect 23436 17106 23492 17500
rect 23436 17054 23438 17106
rect 23490 17054 23492 17106
rect 23436 17042 23492 17054
rect 23660 17220 23716 17230
rect 23660 17106 23716 17164
rect 23660 17054 23662 17106
rect 23714 17054 23716 17106
rect 23660 17042 23716 17054
rect 23772 16996 23828 17006
rect 23772 16902 23828 16940
rect 23996 16884 24052 16894
rect 24220 16884 24276 16894
rect 24052 16828 24164 16884
rect 23996 16818 24052 16828
rect 23548 16772 23604 16782
rect 23548 16678 23604 16716
rect 23100 16146 23156 16156
rect 23996 16212 24052 16222
rect 23996 16118 24052 16156
rect 23212 16098 23268 16110
rect 23212 16046 23214 16098
rect 23266 16046 23268 16098
rect 22092 15428 22148 15438
rect 21980 15426 22148 15428
rect 21980 15374 22094 15426
rect 22146 15374 22148 15426
rect 21980 15372 22148 15374
rect 22092 15362 22148 15372
rect 23212 15316 23268 16046
rect 23212 15250 23268 15260
rect 24108 15204 24164 16828
rect 24220 16790 24276 16828
rect 24332 15316 24388 15326
rect 24668 15316 24724 18286
rect 28140 18338 28196 19068
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 28140 18286 28142 18338
rect 28194 18286 28196 18338
rect 28140 18274 28196 18286
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 24388 15314 24724 15316
rect 24388 15262 24670 15314
rect 24722 15262 24724 15314
rect 24388 15260 24724 15262
rect 24220 15204 24276 15242
rect 24108 15148 24220 15204
rect 24220 15138 24276 15148
rect 22988 14756 23044 14766
rect 22988 14662 23044 14700
rect 21756 13806 21758 13858
rect 21810 13806 21812 13858
rect 21756 13794 21812 13806
rect 23100 14418 23156 14430
rect 23100 14366 23102 14418
rect 23154 14366 23156 14418
rect 21084 13746 21364 13748
rect 21084 13694 21086 13746
rect 21138 13694 21364 13746
rect 21084 13692 21364 13694
rect 21084 13682 21140 13692
rect 23100 13636 23156 14366
rect 24332 13970 24388 15260
rect 24668 15250 24724 15260
rect 26124 16884 26180 16894
rect 26124 16210 26180 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 26124 16158 26126 16210
rect 26178 16158 26180 16210
rect 24332 13918 24334 13970
rect 24386 13918 24388 13970
rect 24332 13906 24388 13918
rect 25228 15204 25284 15214
rect 23100 13570 23156 13580
rect 23884 13636 23940 13646
rect 23884 13542 23940 13580
rect 24556 13636 24612 13646
rect 20748 13076 20804 13086
rect 20524 13074 20804 13076
rect 20524 13022 20750 13074
rect 20802 13022 20804 13074
rect 20524 13020 20804 13022
rect 20748 12740 20804 13020
rect 21308 12740 21364 12750
rect 20748 12738 21364 12740
rect 20748 12686 21310 12738
rect 21362 12686 21364 12738
rect 20748 12684 21364 12686
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 21308 8428 21364 12684
rect 21644 12738 21700 12750
rect 21644 12686 21646 12738
rect 21698 12686 21700 12738
rect 21644 8428 21700 12686
rect 21084 8372 21364 8428
rect 21420 8372 21700 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 21084 4338 21140 8372
rect 21084 4286 21086 4338
rect 21138 4286 21140 4338
rect 21084 4274 21140 4286
rect 20860 4116 20916 4126
rect 19740 3556 19796 3566
rect 19628 3554 19796 3556
rect 19628 3502 19742 3554
rect 19794 3502 19796 3554
rect 19628 3500 19796 3502
rect 19740 3490 19796 3500
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 4060
rect 21420 3554 21476 8372
rect 22092 4116 22148 4126
rect 22092 4022 22148 4060
rect 24220 4116 24276 4126
rect 21420 3502 21422 3554
rect 21474 3502 21476 3554
rect 21420 3490 21476 3502
rect 21532 3668 21588 3678
rect 21532 800 21588 3612
rect 22428 3668 22484 3678
rect 22428 3574 22484 3612
rect 23548 3668 23604 3678
rect 23548 800 23604 3612
rect 24220 800 24276 4060
rect 24556 3554 24612 13580
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24892 5236 24948 5246
rect 24892 800 24948 5180
rect 25228 4338 25284 15148
rect 26124 8428 26180 16158
rect 26572 15874 26628 15886
rect 26572 15822 26574 15874
rect 26626 15822 26628 15874
rect 26460 15316 26516 15326
rect 26572 15316 26628 15822
rect 26516 15260 26628 15316
rect 26460 15250 26516 15260
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 40236 13858 40292 13870
rect 40236 13806 40238 13858
rect 40290 13806 40292 13858
rect 40236 13524 40292 13806
rect 40236 13458 40292 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 25340 8372 26180 8428
rect 25340 5122 25396 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 26124 5236 26180 5246
rect 26124 5142 26180 5180
rect 25340 5070 25342 5122
rect 25394 5070 25396 5122
rect 25340 5058 25396 5070
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 20832 0 20944 800
rect 21504 0 21616 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 24864 0 24976 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 17500 37436 17556 37492
rect 16828 36652 16884 36708
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 14588 28642 14644 28644
rect 14588 28590 14590 28642
rect 14590 28590 14642 28642
rect 14642 28590 14644 28642
rect 14588 28588 14644 28590
rect 4172 28252 4228 28308
rect 1932 25564 1988 25620
rect 2044 24892 2100 24948
rect 16716 28476 16772 28532
rect 17388 28476 17444 28532
rect 17500 28588 17556 28644
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 16828 26908 16884 26964
rect 17388 26908 17444 26964
rect 4284 26290 4340 26292
rect 4284 26238 4286 26290
rect 4286 26238 4338 26290
rect 4338 26238 4340 26290
rect 4284 26236 4340 26238
rect 12684 26236 12740 26292
rect 13580 26124 13636 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 25340 4340 25396
rect 15596 26124 15652 26180
rect 15932 26236 15988 26292
rect 14812 25676 14868 25732
rect 15260 26012 15316 26068
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 12908 22482 12964 22484
rect 12908 22430 12910 22482
rect 12910 22430 12962 22482
rect 12962 22430 12964 22482
rect 12908 22428 12964 22430
rect 14700 24108 14756 24164
rect 10108 21756 10164 21812
rect 11676 21868 11732 21924
rect 10780 21644 10836 21700
rect 11004 21756 11060 21812
rect 14028 22482 14084 22484
rect 14028 22430 14030 22482
rect 14030 22430 14082 22482
rect 14082 22430 14084 22482
rect 14028 22428 14084 22430
rect 14588 22428 14644 22484
rect 14924 22428 14980 22484
rect 14140 22146 14196 22148
rect 14140 22094 14142 22146
rect 14142 22094 14194 22146
rect 14194 22094 14196 22146
rect 14140 22092 14196 22094
rect 13580 21756 13636 21812
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4172 20524 4228 20580
rect 14252 21810 14308 21812
rect 14252 21758 14254 21810
rect 14254 21758 14306 21810
rect 14306 21758 14308 21810
rect 14252 21756 14308 21758
rect 13580 20300 13636 20356
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 1932 18226 1988 18228
rect 1932 18174 1934 18226
rect 1934 18174 1986 18226
rect 1986 18174 1988 18226
rect 1932 18172 1988 18174
rect 11340 18338 11396 18340
rect 11340 18286 11342 18338
rect 11342 18286 11394 18338
rect 11394 18286 11396 18338
rect 11340 18284 11396 18286
rect 13916 19964 13972 20020
rect 13916 19404 13972 19460
rect 14812 20972 14868 21028
rect 16044 26178 16100 26180
rect 16044 26126 16046 26178
rect 16046 26126 16098 26178
rect 16098 26126 16100 26178
rect 16044 26124 16100 26126
rect 16828 26012 16884 26068
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18508 37490 18564 37492
rect 18508 37438 18510 37490
rect 18510 37438 18562 37490
rect 18562 37438 18564 37490
rect 18508 37436 18564 37438
rect 20860 38220 20916 38276
rect 22092 38274 22148 38276
rect 22092 38222 22094 38274
rect 22094 38222 22146 38274
rect 22146 38222 22148 38274
rect 22092 38220 22148 38222
rect 24220 38220 24276 38276
rect 20188 37436 20244 37492
rect 18060 36706 18116 36708
rect 18060 36654 18062 36706
rect 18062 36654 18114 36706
rect 18114 36654 18116 36706
rect 18060 36652 18116 36654
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 17724 28530 17780 28532
rect 17724 28478 17726 28530
rect 17726 28478 17778 28530
rect 17778 28478 17780 28530
rect 17724 28476 17780 28478
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 18508 28642 18564 28644
rect 18508 28590 18510 28642
rect 18510 28590 18562 28642
rect 18562 28590 18564 28642
rect 18508 28588 18564 28590
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17836 27804 17892 27860
rect 18620 27858 18676 27860
rect 18620 27806 18622 27858
rect 18622 27806 18674 27858
rect 18674 27806 18676 27858
rect 18620 27804 18676 27806
rect 21420 37490 21476 37492
rect 21420 37438 21422 37490
rect 21422 37438 21474 37490
rect 21474 37438 21476 37490
rect 21420 37436 21476 37438
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 24892 37436 24948 37492
rect 19292 26796 19348 26852
rect 20524 26796 20580 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19740 26514 19796 26516
rect 19740 26462 19742 26514
rect 19742 26462 19794 26514
rect 19794 26462 19796 26514
rect 19740 26460 19796 26462
rect 21308 27804 21364 27860
rect 20636 26460 20692 26516
rect 17500 26124 17556 26180
rect 16380 25676 16436 25732
rect 16828 25618 16884 25620
rect 16828 25566 16830 25618
rect 16830 25566 16882 25618
rect 16882 25566 16884 25618
rect 16828 25564 16884 25566
rect 17724 26012 17780 26068
rect 17612 25676 17668 25732
rect 16044 25004 16100 25060
rect 16268 24892 16324 24948
rect 16604 24556 16660 24612
rect 16268 24162 16324 24164
rect 16268 24110 16270 24162
rect 16270 24110 16322 24162
rect 16322 24110 16324 24162
rect 16268 24108 16324 24110
rect 15260 22428 15316 22484
rect 15036 22092 15092 22148
rect 15596 22428 15652 22484
rect 16044 22092 16100 22148
rect 15820 21698 15876 21700
rect 15820 21646 15822 21698
rect 15822 21646 15874 21698
rect 15874 21646 15876 21698
rect 15820 21644 15876 21646
rect 15708 21308 15764 21364
rect 15148 20076 15204 20132
rect 15036 19964 15092 20020
rect 15260 20188 15316 20244
rect 18284 25004 18340 25060
rect 17836 24892 17892 24948
rect 17500 24610 17556 24612
rect 17500 24558 17502 24610
rect 17502 24558 17554 24610
rect 17554 24558 17556 24610
rect 17500 24556 17556 24558
rect 17388 23660 17444 23716
rect 17612 23772 17668 23828
rect 17164 23492 17220 23548
rect 16380 23378 16436 23380
rect 16380 23326 16382 23378
rect 16382 23326 16434 23378
rect 16434 23326 16436 23378
rect 16380 23324 16436 23326
rect 16156 20802 16212 20804
rect 16156 20750 16158 20802
rect 16158 20750 16210 20802
rect 16210 20750 16212 20802
rect 16156 20748 16212 20750
rect 15372 19964 15428 20020
rect 15596 20076 15652 20132
rect 15820 19852 15876 19908
rect 15932 20130 15988 20132
rect 15932 20078 15934 20130
rect 15934 20078 15986 20130
rect 15986 20078 15988 20130
rect 15932 20076 15988 20078
rect 14140 18620 14196 18676
rect 14252 18396 14308 18452
rect 13916 18338 13972 18340
rect 13916 18286 13918 18338
rect 13918 18286 13970 18338
rect 13970 18286 13972 18338
rect 13916 18284 13972 18286
rect 13804 18172 13860 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4284 17612 4340 17668
rect 10892 17612 10948 17668
rect 13020 17388 13076 17444
rect 14364 18284 14420 18340
rect 14476 17724 14532 17780
rect 14252 17612 14308 17668
rect 14812 18674 14868 18676
rect 14812 18622 14814 18674
rect 14814 18622 14866 18674
rect 14866 18622 14868 18674
rect 14812 18620 14868 18622
rect 15372 18562 15428 18564
rect 15372 18510 15374 18562
rect 15374 18510 15426 18562
rect 15426 18510 15428 18562
rect 15372 18508 15428 18510
rect 14924 18396 14980 18452
rect 14700 18284 14756 18340
rect 14588 17612 14644 17668
rect 15260 18284 15316 18340
rect 16492 22092 16548 22148
rect 16380 20076 16436 20132
rect 16268 19628 16324 19684
rect 16716 21868 16772 21924
rect 18956 25004 19012 25060
rect 18396 24946 18452 24948
rect 18396 24894 18398 24946
rect 18398 24894 18450 24946
rect 18450 24894 18452 24946
rect 18396 24892 18452 24894
rect 20188 26290 20244 26292
rect 20188 26238 20190 26290
rect 20190 26238 20242 26290
rect 20242 26238 20244 26290
rect 20188 26236 20244 26238
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19068 24892 19124 24948
rect 18732 24780 18788 24836
rect 17836 23548 17892 23604
rect 18060 24722 18116 24724
rect 18060 24670 18062 24722
rect 18062 24670 18114 24722
rect 18114 24670 18116 24722
rect 18060 24668 18116 24670
rect 17612 23324 17668 23380
rect 17388 22146 17444 22148
rect 17388 22094 17390 22146
rect 17390 22094 17442 22146
rect 17442 22094 17444 22146
rect 17388 22092 17444 22094
rect 18060 23660 18116 23716
rect 18620 23826 18676 23828
rect 18620 23774 18622 23826
rect 18622 23774 18674 23826
rect 18674 23774 18676 23826
rect 18620 23772 18676 23774
rect 18508 23324 18564 23380
rect 18620 23548 18676 23604
rect 18844 24668 18900 24724
rect 18956 24556 19012 24612
rect 19740 24108 19796 24164
rect 18060 21756 18116 21812
rect 17836 21586 17892 21588
rect 17836 21534 17838 21586
rect 17838 21534 17890 21586
rect 17890 21534 17892 21586
rect 17836 21532 17892 21534
rect 16716 21308 16772 21364
rect 17500 21362 17556 21364
rect 17500 21310 17502 21362
rect 17502 21310 17554 21362
rect 17554 21310 17556 21362
rect 17500 21308 17556 21310
rect 18732 20636 18788 20692
rect 18844 20972 18900 21028
rect 17948 20524 18004 20580
rect 17724 20130 17780 20132
rect 17724 20078 17726 20130
rect 17726 20078 17778 20130
rect 17778 20078 17780 20130
rect 17724 20076 17780 20078
rect 17388 20018 17444 20020
rect 17388 19966 17390 20018
rect 17390 19966 17442 20018
rect 17442 19966 17444 20018
rect 17388 19964 17444 19966
rect 16044 19404 16100 19460
rect 16828 19628 16884 19684
rect 17388 19404 17444 19460
rect 17276 18508 17332 18564
rect 16268 18226 16324 18228
rect 16268 18174 16270 18226
rect 16270 18174 16322 18226
rect 16322 18174 16324 18226
rect 16268 18172 16324 18174
rect 15260 17666 15316 17668
rect 15260 17614 15262 17666
rect 15262 17614 15314 17666
rect 15314 17614 15316 17666
rect 15260 17612 15316 17614
rect 14476 17554 14532 17556
rect 14476 17502 14478 17554
rect 14478 17502 14530 17554
rect 14530 17502 14532 17554
rect 14476 17500 14532 17502
rect 15148 17442 15204 17444
rect 15148 17390 15150 17442
rect 15150 17390 15202 17442
rect 15202 17390 15204 17442
rect 15148 17388 15204 17390
rect 15708 17666 15764 17668
rect 15708 17614 15710 17666
rect 15710 17614 15762 17666
rect 15762 17614 15764 17666
rect 15708 17612 15764 17614
rect 16156 17666 16212 17668
rect 16156 17614 16158 17666
rect 16158 17614 16210 17666
rect 16210 17614 16212 17666
rect 16156 17612 16212 17614
rect 16492 18060 16548 18116
rect 18060 18956 18116 19012
rect 17724 18562 17780 18564
rect 17724 18510 17726 18562
rect 17726 18510 17778 18562
rect 17778 18510 17780 18562
rect 17724 18508 17780 18510
rect 17276 17724 17332 17780
rect 16604 17612 16660 17668
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 12460 16044 12516 16100
rect 11788 15484 11844 15540
rect 14252 15484 14308 15540
rect 14588 16828 14644 16884
rect 14700 15484 14756 15540
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 15036 15538 15092 15540
rect 15036 15486 15038 15538
rect 15038 15486 15090 15538
rect 15090 15486 15092 15538
rect 15036 15484 15092 15486
rect 17388 17612 17444 17668
rect 17836 17724 17892 17780
rect 16716 16828 16772 16884
rect 17500 16098 17556 16100
rect 17500 16046 17502 16098
rect 17502 16046 17554 16098
rect 17554 16046 17556 16098
rect 17500 16044 17556 16046
rect 18732 20412 18788 20468
rect 18172 18172 18228 18228
rect 18620 20130 18676 20132
rect 18620 20078 18622 20130
rect 18622 20078 18674 20130
rect 18674 20078 18676 20130
rect 18620 20076 18676 20078
rect 18508 19852 18564 19908
rect 18508 18450 18564 18452
rect 18508 18398 18510 18450
rect 18510 18398 18562 18450
rect 18562 18398 18564 18450
rect 18508 18396 18564 18398
rect 18284 17724 18340 17780
rect 18620 17666 18676 17668
rect 18620 17614 18622 17666
rect 18622 17614 18674 17666
rect 18674 17614 18676 17666
rect 18620 17612 18676 17614
rect 24668 28476 24724 28532
rect 21756 27858 21812 27860
rect 21756 27806 21758 27858
rect 21758 27806 21810 27858
rect 21810 27806 21812 27858
rect 21756 27804 21812 27806
rect 22316 27804 22372 27860
rect 22540 27746 22596 27748
rect 22540 27694 22542 27746
rect 22542 27694 22594 27746
rect 22594 27694 22596 27746
rect 22540 27692 22596 27694
rect 21532 26962 21588 26964
rect 21532 26910 21534 26962
rect 21534 26910 21586 26962
rect 21586 26910 21588 26962
rect 21532 26908 21588 26910
rect 22316 26796 22372 26852
rect 23548 26908 23604 26964
rect 20636 26290 20692 26292
rect 20636 26238 20638 26290
rect 20638 26238 20690 26290
rect 20690 26238 20692 26290
rect 20636 26236 20692 26238
rect 20412 24108 20468 24164
rect 20748 23772 20804 23828
rect 21308 26236 21364 26292
rect 21196 24780 21252 24836
rect 23436 26514 23492 26516
rect 23436 26462 23438 26514
rect 23438 26462 23490 26514
rect 23490 26462 23492 26514
rect 23436 26460 23492 26462
rect 24332 26908 24388 26964
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 26236 37884 26292 37940
rect 27468 37938 27524 37940
rect 27468 37886 27470 37938
rect 27470 37886 27522 37938
rect 27522 37886 27524 37938
rect 27468 37884 27524 37886
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 25228 28476 25284 28532
rect 24556 27020 24612 27076
rect 25116 26460 25172 26516
rect 25452 27692 25508 27748
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 25564 26962 25620 26964
rect 25564 26910 25566 26962
rect 25566 26910 25618 26962
rect 25618 26910 25620 26962
rect 25564 26908 25620 26910
rect 25340 26796 25396 26852
rect 23212 26290 23268 26292
rect 23212 26238 23214 26290
rect 23214 26238 23266 26290
rect 23266 26238 23268 26290
rect 23212 26236 23268 26238
rect 23212 25228 23268 25284
rect 21420 24892 21476 24948
rect 20076 23660 20132 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19180 20748 19236 20804
rect 18844 20188 18900 20244
rect 19292 20412 19348 20468
rect 19852 23154 19908 23156
rect 19852 23102 19854 23154
rect 19854 23102 19906 23154
rect 19906 23102 19908 23154
rect 19852 23100 19908 23102
rect 20412 22988 20468 23044
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19852 21756 19908 21812
rect 19628 21308 19684 21364
rect 19852 20972 19908 21028
rect 20300 21474 20356 21476
rect 20300 21422 20302 21474
rect 20302 21422 20354 21474
rect 20354 21422 20356 21474
rect 20300 21420 20356 21422
rect 20188 20802 20244 20804
rect 20188 20750 20190 20802
rect 20190 20750 20242 20802
rect 20242 20750 20244 20802
rect 20188 20748 20244 20750
rect 20076 20690 20132 20692
rect 20076 20638 20078 20690
rect 20078 20638 20130 20690
rect 20130 20638 20132 20690
rect 20076 20636 20132 20638
rect 19964 20578 20020 20580
rect 19964 20526 19966 20578
rect 19966 20526 20018 20578
rect 20018 20526 20020 20578
rect 19964 20524 20020 20526
rect 19516 20412 19572 20468
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20636 20972 20692 21028
rect 19964 20242 20020 20244
rect 19964 20190 19966 20242
rect 19966 20190 20018 20242
rect 20018 20190 20020 20242
rect 19964 20188 20020 20190
rect 19404 20130 19460 20132
rect 19404 20078 19406 20130
rect 19406 20078 19458 20130
rect 19458 20078 19460 20130
rect 19404 20076 19460 20078
rect 19404 19740 19460 19796
rect 19292 19292 19348 19348
rect 19628 19964 19684 20020
rect 18844 18284 18900 18340
rect 20076 20018 20132 20020
rect 20076 19966 20078 20018
rect 20078 19966 20130 20018
rect 20130 19966 20132 20018
rect 20076 19964 20132 19966
rect 21084 23154 21140 23156
rect 21084 23102 21086 23154
rect 21086 23102 21138 23154
rect 21138 23102 21140 23154
rect 21084 23100 21140 23102
rect 20972 20748 21028 20804
rect 22540 24946 22596 24948
rect 22540 24894 22542 24946
rect 22542 24894 22594 24946
rect 22594 24894 22596 24946
rect 22540 24892 22596 24894
rect 22316 24834 22372 24836
rect 22316 24782 22318 24834
rect 22318 24782 22370 24834
rect 22370 24782 22372 24834
rect 22316 24780 22372 24782
rect 22204 24556 22260 24612
rect 22204 23714 22260 23716
rect 22204 23662 22206 23714
rect 22206 23662 22258 23714
rect 22258 23662 22260 23714
rect 22204 23660 22260 23662
rect 22428 23212 22484 23268
rect 21868 21756 21924 21812
rect 21532 21532 21588 21588
rect 21532 20412 21588 20468
rect 21644 20972 21700 21028
rect 20412 19852 20468 19908
rect 20188 19292 20244 19348
rect 19740 18956 19796 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 18060 16322 18116 16324
rect 18060 16270 18062 16322
rect 18062 16270 18114 16322
rect 18114 16270 18116 16322
rect 18060 16268 18116 16270
rect 18396 15932 18452 15988
rect 17276 15820 17332 15876
rect 17388 15372 17444 15428
rect 16604 15314 16660 15316
rect 16604 15262 16606 15314
rect 16606 15262 16658 15314
rect 16658 15262 16660 15314
rect 16604 15260 16660 15262
rect 16716 15202 16772 15204
rect 16716 15150 16718 15202
rect 16718 15150 16770 15202
rect 16770 15150 16772 15202
rect 16716 15148 16772 15150
rect 17500 15260 17556 15316
rect 18284 15708 18340 15764
rect 18732 15820 18788 15876
rect 18956 17778 19012 17780
rect 18956 17726 18958 17778
rect 18958 17726 19010 17778
rect 19010 17726 19012 17778
rect 18956 17724 19012 17726
rect 18732 15372 18788 15428
rect 14700 14530 14756 14532
rect 14700 14478 14702 14530
rect 14702 14478 14754 14530
rect 14754 14478 14756 14530
rect 14700 14476 14756 14478
rect 16380 14476 16436 14532
rect 16828 13970 16884 13972
rect 16828 13918 16830 13970
rect 16830 13918 16882 13970
rect 16882 13918 16884 13970
rect 16828 13916 16884 13918
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 17948 14530 18004 14532
rect 17948 14478 17950 14530
rect 17950 14478 18002 14530
rect 18002 14478 18004 14530
rect 17948 14476 18004 14478
rect 17500 13916 17556 13972
rect 18508 15314 18564 15316
rect 18508 15262 18510 15314
rect 18510 15262 18562 15314
rect 18562 15262 18564 15314
rect 18508 15260 18564 15262
rect 18620 15202 18676 15204
rect 18620 15150 18622 15202
rect 18622 15150 18674 15202
rect 18674 15150 18676 15202
rect 18620 15148 18676 15150
rect 20188 18620 20244 18676
rect 20412 19180 20468 19236
rect 20300 18450 20356 18452
rect 20300 18398 20302 18450
rect 20302 18398 20354 18450
rect 20354 18398 20356 18450
rect 20300 18396 20356 18398
rect 19516 17442 19572 17444
rect 19516 17390 19518 17442
rect 19518 17390 19570 17442
rect 19570 17390 19572 17442
rect 19516 17388 19572 17390
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20076 17052 20132 17108
rect 19292 16828 19348 16884
rect 19180 15986 19236 15988
rect 19180 15934 19182 15986
rect 19182 15934 19234 15986
rect 19234 15934 19236 15986
rect 19180 15932 19236 15934
rect 19404 16098 19460 16100
rect 19404 16046 19406 16098
rect 19406 16046 19458 16098
rect 19458 16046 19460 16098
rect 19404 16044 19460 16046
rect 19404 15820 19460 15876
rect 21420 20018 21476 20020
rect 21420 19966 21422 20018
rect 21422 19966 21474 20018
rect 21474 19966 21476 20018
rect 21420 19964 21476 19966
rect 21532 19740 21588 19796
rect 20636 18284 20692 18340
rect 20972 18620 21028 18676
rect 24108 25228 24164 25284
rect 23772 24892 23828 24948
rect 22540 21756 22596 21812
rect 21980 21420 22036 21476
rect 23548 23324 23604 23380
rect 23212 23212 23268 23268
rect 26012 26850 26068 26852
rect 26012 26798 26014 26850
rect 26014 26798 26066 26850
rect 26066 26798 26068 26850
rect 26012 26796 26068 26798
rect 27244 26124 27300 26180
rect 28364 26178 28420 26180
rect 28364 26126 28366 26178
rect 28366 26126 28418 26178
rect 28418 26126 28420 26178
rect 28364 26124 28420 26126
rect 40012 26236 40068 26292
rect 37660 26124 37716 26180
rect 27356 26012 27412 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 24220 24556 24276 24612
rect 25900 24892 25956 24948
rect 26124 25282 26180 25284
rect 26124 25230 26126 25282
rect 26126 25230 26178 25282
rect 26178 25230 26180 25282
rect 26124 25228 26180 25230
rect 22876 20972 22932 21028
rect 22204 20860 22260 20916
rect 22316 20636 22372 20692
rect 21868 20412 21924 20468
rect 21756 20300 21812 20356
rect 21084 18562 21140 18564
rect 21084 18510 21086 18562
rect 21086 18510 21138 18562
rect 21138 18510 21140 18562
rect 21084 18508 21140 18510
rect 20972 18396 21028 18452
rect 21980 20130 22036 20132
rect 21980 20078 21982 20130
rect 21982 20078 22034 20130
rect 22034 20078 22036 20130
rect 21980 20076 22036 20078
rect 22540 20578 22596 20580
rect 22540 20526 22542 20578
rect 22542 20526 22594 20578
rect 22594 20526 22596 20578
rect 22540 20524 22596 20526
rect 22092 19964 22148 20020
rect 22876 20188 22932 20244
rect 23660 20188 23716 20244
rect 21868 19234 21924 19236
rect 21868 19182 21870 19234
rect 21870 19182 21922 19234
rect 21922 19182 21924 19234
rect 21868 19180 21924 19182
rect 21644 18284 21700 18340
rect 22540 19010 22596 19012
rect 22540 18958 22542 19010
rect 22542 18958 22594 19010
rect 22594 18958 22596 19010
rect 22540 18956 22596 18958
rect 20524 17052 20580 17108
rect 22204 17500 22260 17556
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19964 15484 20020 15540
rect 19516 15260 19572 15316
rect 19628 14306 19684 14308
rect 19628 14254 19630 14306
rect 19630 14254 19682 14306
rect 19682 14254 19684 14306
rect 19628 14252 19684 14254
rect 20300 15314 20356 15316
rect 20300 15262 20302 15314
rect 20302 15262 20354 15314
rect 20354 15262 20356 15314
rect 20300 15260 20356 15262
rect 21532 17388 21588 17444
rect 20748 17276 20804 17332
rect 21196 17106 21252 17108
rect 21196 17054 21198 17106
rect 21198 17054 21250 17106
rect 21250 17054 21252 17106
rect 21196 17052 21252 17054
rect 21420 17106 21476 17108
rect 21420 17054 21422 17106
rect 21422 17054 21474 17106
rect 21474 17054 21476 17106
rect 21420 17052 21476 17054
rect 22316 17388 22372 17444
rect 24444 23042 24500 23044
rect 24444 22990 24446 23042
rect 24446 22990 24498 23042
rect 24498 22990 24500 23042
rect 24444 22988 24500 22990
rect 24444 22204 24500 22260
rect 27356 23996 27412 24052
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 28588 24050 28644 24052
rect 28588 23998 28590 24050
rect 28590 23998 28642 24050
rect 28642 23998 28644 24050
rect 28588 23996 28644 23998
rect 40012 24220 40068 24276
rect 37660 23996 37716 24052
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 25340 22204 25396 22260
rect 25788 22258 25844 22260
rect 25788 22206 25790 22258
rect 25790 22206 25842 22258
rect 25842 22206 25844 22258
rect 25788 22204 25844 22206
rect 24108 21810 24164 21812
rect 24108 21758 24110 21810
rect 24110 21758 24162 21810
rect 24162 21758 24164 21810
rect 24108 21756 24164 21758
rect 23884 20524 23940 20580
rect 24332 21196 24388 21252
rect 24108 20188 24164 20244
rect 24332 20860 24388 20916
rect 25228 20860 25284 20916
rect 25788 21196 25844 21252
rect 24668 20130 24724 20132
rect 24668 20078 24670 20130
rect 24670 20078 24722 20130
rect 24722 20078 24724 20130
rect 24668 20076 24724 20078
rect 24556 19740 24612 19796
rect 26348 20690 26404 20692
rect 26348 20638 26350 20690
rect 26350 20638 26402 20690
rect 26402 20638 26404 20690
rect 26348 20636 26404 20638
rect 25340 20130 25396 20132
rect 25340 20078 25342 20130
rect 25342 20078 25394 20130
rect 25394 20078 25396 20130
rect 25340 20076 25396 20078
rect 24780 19068 24836 19124
rect 22652 18396 22708 18452
rect 22428 17276 22484 17332
rect 22540 18284 22596 18340
rect 22540 17164 22596 17220
rect 23660 18396 23716 18452
rect 24220 19010 24276 19012
rect 24220 18958 24222 19010
rect 24222 18958 24274 19010
rect 24274 18958 24276 19010
rect 24220 18956 24276 18958
rect 23996 17836 24052 17892
rect 24668 18396 24724 18452
rect 25788 19292 25844 19348
rect 25900 19122 25956 19124
rect 25900 19070 25902 19122
rect 25902 19070 25954 19122
rect 25954 19070 25956 19122
rect 25900 19068 25956 19070
rect 25564 18956 25620 19012
rect 25340 18450 25396 18452
rect 25340 18398 25342 18450
rect 25342 18398 25394 18450
rect 25394 18398 25396 18450
rect 25340 18396 25396 18398
rect 26684 20300 26740 20356
rect 26124 20130 26180 20132
rect 26124 20078 26126 20130
rect 26126 20078 26178 20130
rect 26178 20078 26180 20130
rect 26124 20076 26180 20078
rect 26348 20188 26404 20244
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 27356 21420 27412 21476
rect 28700 21474 28756 21476
rect 28700 21422 28702 21474
rect 28702 21422 28754 21474
rect 28754 21422 28756 21474
rect 28700 21420 28756 21422
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 40012 22204 40068 22260
rect 40012 21532 40068 21588
rect 37884 20972 37940 21028
rect 27356 20914 27412 20916
rect 27356 20862 27358 20914
rect 27358 20862 27410 20914
rect 27410 20862 27412 20914
rect 27356 20860 27412 20862
rect 27132 20188 27188 20244
rect 26236 19794 26292 19796
rect 26236 19742 26238 19794
rect 26238 19742 26290 19794
rect 26290 19742 26292 19794
rect 26236 19740 26292 19742
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 37660 19404 37716 19460
rect 26572 19292 26628 19348
rect 28028 19346 28084 19348
rect 28028 19294 28030 19346
rect 28030 19294 28082 19346
rect 28082 19294 28084 19346
rect 28028 19292 28084 19294
rect 37660 19234 37716 19236
rect 37660 19182 37662 19234
rect 37662 19182 37714 19234
rect 37714 19182 37716 19234
rect 37660 19180 37716 19182
rect 28140 19068 28196 19124
rect 22652 16994 22708 16996
rect 22652 16942 22654 16994
rect 22654 16942 22706 16994
rect 22706 16942 22708 16994
rect 22652 16940 22708 16942
rect 22316 16882 22372 16884
rect 22316 16830 22318 16882
rect 22318 16830 22370 16882
rect 22370 16830 22372 16882
rect 22316 16828 22372 16830
rect 21644 16716 21700 16772
rect 21420 15932 21476 15988
rect 20972 14700 21028 14756
rect 21308 15314 21364 15316
rect 21308 15262 21310 15314
rect 21310 15262 21362 15314
rect 21362 15262 21364 15314
rect 21308 15260 21364 15262
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20412 14306 20468 14308
rect 20412 14254 20414 14306
rect 20414 14254 20466 14306
rect 20466 14254 20468 14306
rect 20412 14252 20468 14254
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 17500 4060 17556 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 18732 4114 18788 4116
rect 18732 4062 18734 4114
rect 18734 4062 18786 4114
rect 18786 4062 18788 4114
rect 18732 4060 18788 4062
rect 22428 16770 22484 16772
rect 22428 16718 22430 16770
rect 22430 16718 22482 16770
rect 22482 16718 22484 16770
rect 22428 16716 22484 16718
rect 23436 17500 23492 17556
rect 22876 17052 22932 17108
rect 23100 17276 23156 17332
rect 22988 16882 23044 16884
rect 22988 16830 22990 16882
rect 22990 16830 23042 16882
rect 23042 16830 23044 16882
rect 22988 16828 23044 16830
rect 22764 16716 22820 16772
rect 23660 17164 23716 17220
rect 23772 16994 23828 16996
rect 23772 16942 23774 16994
rect 23774 16942 23826 16994
rect 23826 16942 23828 16994
rect 23772 16940 23828 16942
rect 23996 16828 24052 16884
rect 23548 16770 23604 16772
rect 23548 16718 23550 16770
rect 23550 16718 23602 16770
rect 23602 16718 23604 16770
rect 23548 16716 23604 16718
rect 23100 16156 23156 16212
rect 23996 16210 24052 16212
rect 23996 16158 23998 16210
rect 23998 16158 24050 16210
rect 24050 16158 24052 16210
rect 23996 16156 24052 16158
rect 23212 15260 23268 15316
rect 24220 16882 24276 16884
rect 24220 16830 24222 16882
rect 24222 16830 24274 16882
rect 24274 16830 24276 16882
rect 24220 16828 24276 16830
rect 40012 18844 40068 18900
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 24332 15260 24388 15316
rect 24220 15202 24276 15204
rect 24220 15150 24222 15202
rect 24222 15150 24274 15202
rect 24274 15150 24276 15202
rect 24220 15148 24276 15150
rect 22988 14754 23044 14756
rect 22988 14702 22990 14754
rect 22990 14702 23042 14754
rect 23042 14702 23044 14754
rect 22988 14700 23044 14702
rect 26124 16828 26180 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 25228 15148 25284 15204
rect 23100 13580 23156 13636
rect 23884 13634 23940 13636
rect 23884 13582 23886 13634
rect 23886 13582 23938 13634
rect 23938 13582 23940 13634
rect 23884 13580 23940 13582
rect 24556 13580 24612 13636
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20860 4060 20916 4116
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22092 4114 22148 4116
rect 22092 4062 22094 4114
rect 22094 4062 22146 4114
rect 22146 4062 22148 4114
rect 22092 4060 22148 4062
rect 24220 4060 24276 4116
rect 21532 3612 21588 3668
rect 22428 3666 22484 3668
rect 22428 3614 22430 3666
rect 22430 3614 22482 3666
rect 22482 3614 22484 3666
rect 22428 3612 22484 3614
rect 23548 3612 23604 3668
rect 24892 5180 24948 5236
rect 26460 15260 26516 15316
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 40236 13468 40292 13524
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26124 5234 26180 5236
rect 26124 5182 26126 5234
rect 26126 5182 26178 5234
rect 26178 5182 26180 5234
rect 26124 5180 26180 5182
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 20850 38220 20860 38276
rect 20916 38220 22092 38276
rect 22148 38220 22158 38276
rect 24210 38220 24220 38276
rect 24276 38220 25564 38276
rect 25620 38220 25630 38276
rect 26226 37884 26236 37940
rect 26292 37884 27468 37940
rect 27524 37884 27534 37940
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 17490 37436 17500 37492
rect 17556 37436 18508 37492
rect 18564 37436 18574 37492
rect 20178 37436 20188 37492
rect 20244 37436 21420 37492
rect 21476 37436 21486 37492
rect 24882 37436 24892 37492
rect 24948 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 16818 36652 16828 36708
rect 16884 36652 18060 36708
rect 18116 36652 18126 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 14578 28588 14588 28644
rect 14644 28588 17500 28644
rect 17556 28588 18508 28644
rect 18564 28588 18574 28644
rect 16706 28476 16716 28532
rect 16772 28476 17388 28532
rect 17444 28476 17724 28532
rect 17780 28476 17790 28532
rect 24658 28476 24668 28532
rect 24724 28476 25228 28532
rect 25284 28476 25294 28532
rect 0 28308 800 28336
rect 0 28252 4172 28308
rect 4228 28252 4238 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 17826 27804 17836 27860
rect 17892 27804 18620 27860
rect 18676 27804 21308 27860
rect 21364 27804 21756 27860
rect 21812 27804 22316 27860
rect 22372 27804 22382 27860
rect 22530 27692 22540 27748
rect 22596 27692 25452 27748
rect 25508 27692 25518 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 23548 27020 24556 27076
rect 24612 27020 24622 27076
rect 23548 26964 23604 27020
rect 16818 26908 16828 26964
rect 16884 26908 17388 26964
rect 17444 26908 21532 26964
rect 21588 26908 23548 26964
rect 23604 26908 23614 26964
rect 24322 26908 24332 26964
rect 24388 26908 25564 26964
rect 25620 26908 25630 26964
rect 19282 26796 19292 26852
rect 19348 26796 20524 26852
rect 20580 26796 20590 26852
rect 22306 26796 22316 26852
rect 22372 26796 25340 26852
rect 25396 26796 26012 26852
rect 26068 26796 26078 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 19730 26460 19740 26516
rect 19796 26460 20636 26516
rect 20692 26460 20702 26516
rect 23426 26460 23436 26516
rect 23492 26460 25116 26516
rect 25172 26460 25182 26516
rect 41200 26292 42000 26320
rect 4274 26236 4284 26292
rect 4340 26236 12684 26292
rect 12740 26236 15932 26292
rect 15988 26236 15998 26292
rect 20178 26236 20188 26292
rect 20244 26236 20636 26292
rect 20692 26236 20702 26292
rect 21298 26236 21308 26292
rect 21364 26236 23212 26292
rect 23268 26236 23278 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 41200 26208 42000 26236
rect 13570 26124 13580 26180
rect 13636 26124 15596 26180
rect 15652 26124 16044 26180
rect 16100 26124 17500 26180
rect 17556 26124 17566 26180
rect 27234 26124 27244 26180
rect 27300 26124 28364 26180
rect 28420 26124 37660 26180
rect 37716 26124 37726 26180
rect 15250 26012 15260 26068
rect 15316 26012 16828 26068
rect 16884 26012 17724 26068
rect 17780 26012 27356 26068
rect 27412 26012 27422 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14802 25676 14812 25732
rect 14868 25676 15148 25732
rect 16370 25676 16380 25732
rect 16436 25676 17612 25732
rect 17668 25676 17678 25732
rect 0 25620 800 25648
rect 15092 25620 15148 25676
rect 0 25564 1932 25620
rect 1988 25564 1998 25620
rect 15092 25564 16828 25620
rect 16884 25564 16894 25620
rect 0 25536 800 25564
rect 17052 25396 17108 25676
rect 4274 25340 4284 25396
rect 4340 25340 17108 25396
rect 23202 25228 23212 25284
rect 23268 25228 24108 25284
rect 24164 25228 26124 25284
rect 26180 25228 26190 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 16034 25004 16044 25060
rect 16100 25004 18284 25060
rect 18340 25004 18350 25060
rect 18946 25004 18956 25060
rect 19012 25004 19684 25060
rect 0 24948 800 24976
rect 19628 24948 19684 25004
rect 0 24892 2044 24948
rect 2100 24892 2110 24948
rect 16258 24892 16268 24948
rect 16324 24892 17836 24948
rect 17892 24892 18396 24948
rect 18452 24892 19068 24948
rect 19124 24892 19134 24948
rect 19628 24892 21420 24948
rect 21476 24892 21486 24948
rect 22530 24892 22540 24948
rect 22596 24892 23772 24948
rect 23828 24892 25900 24948
rect 25956 24892 25966 24948
rect 0 24864 800 24892
rect 18722 24780 18732 24836
rect 18788 24780 21196 24836
rect 21252 24780 22316 24836
rect 22372 24780 22382 24836
rect 18050 24668 18060 24724
rect 18116 24668 18844 24724
rect 18900 24668 18910 24724
rect 16594 24556 16604 24612
rect 16660 24556 17500 24612
rect 17556 24556 17566 24612
rect 18946 24556 18956 24612
rect 19012 24556 22204 24612
rect 22260 24556 24220 24612
rect 24276 24556 24286 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 41200 24276 42000 24304
rect 40002 24220 40012 24276
rect 40068 24220 42000 24276
rect 41200 24192 42000 24220
rect 14690 24108 14700 24164
rect 14756 24108 16268 24164
rect 16324 24108 16334 24164
rect 19730 24108 19740 24164
rect 19796 24108 20412 24164
rect 20468 24108 20478 24164
rect 27346 23996 27356 24052
rect 27412 23996 28588 24052
rect 28644 23996 37660 24052
rect 37716 23996 37726 24052
rect 17602 23772 17612 23828
rect 17668 23772 18620 23828
rect 18676 23772 18686 23828
rect 19852 23772 20748 23828
rect 20804 23772 20814 23828
rect 19852 23716 19908 23772
rect 17378 23660 17388 23716
rect 17444 23660 18060 23716
rect 18116 23660 19908 23716
rect 20066 23660 20076 23716
rect 20132 23660 22204 23716
rect 22260 23660 22270 23716
rect 17826 23548 17836 23604
rect 17892 23548 18620 23604
rect 18676 23548 18686 23604
rect 17154 23492 17164 23548
rect 17220 23492 17230 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 17164 23436 19404 23492
rect 19460 23436 19470 23492
rect 16370 23324 16380 23380
rect 16436 23324 17612 23380
rect 17668 23324 17678 23380
rect 18498 23324 18508 23380
rect 18564 23324 23548 23380
rect 23604 23324 23614 23380
rect 22418 23212 22428 23268
rect 22484 23212 23212 23268
rect 23268 23212 31948 23268
rect 31892 23156 31948 23212
rect 19842 23100 19852 23156
rect 19908 23100 21084 23156
rect 21140 23100 21150 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 20402 22988 20412 23044
rect 20468 22988 24444 23044
rect 24500 22988 24510 23044
rect 41200 22932 42000 22960
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 12898 22428 12908 22484
rect 12964 22428 14028 22484
rect 14084 22428 14588 22484
rect 14644 22428 14654 22484
rect 14914 22428 14924 22484
rect 14980 22428 15260 22484
rect 15316 22428 15596 22484
rect 15652 22428 15662 22484
rect 41200 22260 42000 22288
rect 24434 22204 24444 22260
rect 24500 22204 25340 22260
rect 25396 22204 25788 22260
rect 25844 22204 25854 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 14130 22092 14140 22148
rect 14196 22092 15036 22148
rect 15092 22092 16044 22148
rect 16100 22092 16110 22148
rect 16482 22092 16492 22148
rect 16548 22092 17388 22148
rect 17444 22092 17454 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 11666 21868 11676 21924
rect 11732 21868 16716 21924
rect 16772 21868 16782 21924
rect 10098 21756 10108 21812
rect 10164 21756 11004 21812
rect 11060 21756 13580 21812
rect 13636 21756 14252 21812
rect 14308 21756 14318 21812
rect 18050 21756 18060 21812
rect 18116 21756 19852 21812
rect 19908 21756 19918 21812
rect 21858 21756 21868 21812
rect 21924 21756 22540 21812
rect 22596 21756 24108 21812
rect 24164 21756 24174 21812
rect 10770 21644 10780 21700
rect 10836 21644 15820 21700
rect 15876 21644 15886 21700
rect 41200 21588 42000 21616
rect 17826 21532 17836 21588
rect 17892 21532 21532 21588
rect 21588 21532 21598 21588
rect 31892 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 31892 21476 31948 21532
rect 41200 21504 42000 21532
rect 20290 21420 20300 21476
rect 20356 21420 21980 21476
rect 22036 21420 22046 21476
rect 27346 21420 27356 21476
rect 27412 21420 28700 21476
rect 28756 21420 31948 21476
rect 15698 21308 15708 21364
rect 15764 21308 16716 21364
rect 16772 21308 17500 21364
rect 17556 21308 19628 21364
rect 19684 21308 19694 21364
rect 24322 21196 24332 21252
rect 24388 21196 25788 21252
rect 25844 21196 25854 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 25788 21028 25844 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 14802 20972 14812 21028
rect 14868 20972 18844 21028
rect 18900 20972 18910 21028
rect 19842 20972 19852 21028
rect 19908 20972 20636 21028
rect 20692 20972 20702 21028
rect 21634 20972 21644 21028
rect 21700 20972 22876 21028
rect 22932 20972 22942 21028
rect 25788 20972 37884 21028
rect 37940 20972 37950 21028
rect 16156 20860 22204 20916
rect 22260 20860 24332 20916
rect 24388 20860 24398 20916
rect 25218 20860 25228 20916
rect 25284 20860 27356 20916
rect 27412 20860 27422 20916
rect 16156 20804 16212 20860
rect 16146 20748 16156 20804
rect 16212 20748 16222 20804
rect 19170 20748 19180 20804
rect 19236 20748 20188 20804
rect 20244 20748 20972 20804
rect 21028 20748 21038 20804
rect 18722 20636 18732 20692
rect 18788 20636 20076 20692
rect 20132 20636 20142 20692
rect 22306 20636 22316 20692
rect 22372 20636 26348 20692
rect 26404 20636 26414 20692
rect 4162 20524 4172 20580
rect 4228 20524 17948 20580
rect 18004 20524 18014 20580
rect 19954 20524 19964 20580
rect 20020 20524 20244 20580
rect 22530 20524 22540 20580
rect 22596 20524 23884 20580
rect 23940 20524 23950 20580
rect 18722 20412 18732 20468
rect 18788 20412 19292 20468
rect 19348 20412 19358 20468
rect 19478 20412 19516 20468
rect 19572 20412 19582 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 13570 20300 13580 20356
rect 13636 20300 15148 20356
rect 15092 20244 15148 20300
rect 15092 20188 15260 20244
rect 15316 20188 15326 20244
rect 18834 20188 18844 20244
rect 18900 20188 19964 20244
rect 20020 20188 20030 20244
rect 20188 20132 20244 20524
rect 21522 20412 21532 20468
rect 21588 20412 21868 20468
rect 21924 20412 21934 20468
rect 21746 20300 21756 20356
rect 21812 20300 26684 20356
rect 26740 20300 26750 20356
rect 22866 20188 22876 20244
rect 22932 20188 23660 20244
rect 23716 20188 23726 20244
rect 24098 20188 24108 20244
rect 24164 20188 26348 20244
rect 26404 20188 27132 20244
rect 27188 20188 27198 20244
rect 15138 20076 15148 20132
rect 15204 20076 15596 20132
rect 15652 20076 15662 20132
rect 15922 20076 15932 20132
rect 15988 20076 16380 20132
rect 16436 20076 16446 20132
rect 17714 20076 17724 20132
rect 17780 20076 18620 20132
rect 18676 20076 18686 20132
rect 19366 20076 19404 20132
rect 19460 20076 19470 20132
rect 20188 20076 21980 20132
rect 22036 20076 22046 20132
rect 24658 20076 24668 20132
rect 24724 20076 25340 20132
rect 25396 20076 26124 20132
rect 26180 20076 26190 20132
rect 18620 20020 18676 20076
rect 13906 19964 13916 20020
rect 13972 19964 15036 20020
rect 15092 19964 15372 20020
rect 15428 19964 17388 20020
rect 17444 19964 17454 20020
rect 18620 19964 19628 20020
rect 19684 19964 20076 20020
rect 20132 19964 20142 20020
rect 21410 19964 21420 20020
rect 21476 19964 22092 20020
rect 22148 19964 22158 20020
rect 15810 19852 15820 19908
rect 15876 19852 18508 19908
rect 18564 19852 19516 19908
rect 19572 19852 20412 19908
rect 20468 19852 20478 19908
rect 19394 19740 19404 19796
rect 19460 19740 21532 19796
rect 21588 19740 21598 19796
rect 24546 19740 24556 19796
rect 24612 19740 26236 19796
rect 26292 19740 26302 19796
rect 16258 19628 16268 19684
rect 16324 19628 16828 19684
rect 16884 19628 16894 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 13906 19404 13916 19460
rect 13972 19404 16044 19460
rect 16100 19404 17388 19460
rect 17444 19404 17454 19460
rect 31892 19404 37660 19460
rect 37716 19404 37726 19460
rect 31892 19348 31948 19404
rect 19282 19292 19292 19348
rect 19348 19292 20188 19348
rect 20244 19292 20254 19348
rect 25778 19292 25788 19348
rect 25844 19292 25854 19348
rect 26562 19292 26572 19348
rect 26628 19292 28028 19348
rect 28084 19292 31948 19348
rect 25788 19236 25844 19292
rect 20402 19180 20412 19236
rect 20468 19180 21868 19236
rect 21924 19180 21934 19236
rect 25788 19180 26908 19236
rect 26852 19124 26908 19180
rect 31892 19180 37660 19236
rect 37716 19180 37726 19236
rect 31892 19124 31948 19180
rect 24770 19068 24780 19124
rect 24836 19068 25900 19124
rect 25956 19068 25966 19124
rect 26852 19068 28140 19124
rect 28196 19068 31948 19124
rect 18050 18956 18060 19012
rect 18116 18956 19740 19012
rect 19796 18956 19806 19012
rect 22530 18956 22540 19012
rect 22596 18956 24220 19012
rect 24276 18956 25564 19012
rect 25620 18956 25630 19012
rect 41200 18900 42000 18928
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 14130 18620 14140 18676
rect 14196 18620 14812 18676
rect 14868 18620 14878 18676
rect 20178 18620 20188 18676
rect 20244 18620 20972 18676
rect 21028 18620 21038 18676
rect 15362 18508 15372 18564
rect 15428 18508 17276 18564
rect 17332 18508 17342 18564
rect 17714 18508 17724 18564
rect 17780 18508 21084 18564
rect 21140 18508 21150 18564
rect 14242 18396 14252 18452
rect 14308 18396 14924 18452
rect 14980 18396 14990 18452
rect 18498 18396 18508 18452
rect 18564 18396 20300 18452
rect 20356 18396 20366 18452
rect 20962 18396 20972 18452
rect 21028 18396 22652 18452
rect 22708 18396 22718 18452
rect 23650 18396 23660 18452
rect 23716 18396 24668 18452
rect 24724 18396 25340 18452
rect 25396 18396 25406 18452
rect 11330 18284 11340 18340
rect 11396 18284 13916 18340
rect 13972 18284 14364 18340
rect 14420 18284 14430 18340
rect 14690 18284 14700 18340
rect 14756 18284 15260 18340
rect 15316 18284 18844 18340
rect 18900 18284 18910 18340
rect 20626 18284 20636 18340
rect 20692 18284 21644 18340
rect 21700 18284 22540 18340
rect 22596 18284 22606 18340
rect 0 18228 800 18256
rect 0 18172 1932 18228
rect 1988 18172 1998 18228
rect 13794 18172 13804 18228
rect 13860 18172 16268 18228
rect 16324 18172 18172 18228
rect 18228 18172 18238 18228
rect 0 18144 800 18172
rect 16492 18116 16548 18172
rect 16482 18060 16492 18116
rect 16548 18060 16558 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 15932 17836 23996 17892
rect 24052 17836 24062 17892
rect 15932 17780 15988 17836
rect 14466 17724 14476 17780
rect 14532 17724 15988 17780
rect 17266 17724 17276 17780
rect 17332 17724 17836 17780
rect 17892 17724 18284 17780
rect 18340 17724 18956 17780
rect 19012 17724 19022 17780
rect 15932 17668 15988 17724
rect 4274 17612 4284 17668
rect 4340 17612 10892 17668
rect 10948 17612 14252 17668
rect 14308 17612 14318 17668
rect 14578 17612 14588 17668
rect 14644 17612 15260 17668
rect 15316 17612 15326 17668
rect 15698 17612 15708 17668
rect 15764 17612 15988 17668
rect 16146 17612 16156 17668
rect 16212 17612 16222 17668
rect 16594 17612 16604 17668
rect 16660 17612 17388 17668
rect 17444 17612 18620 17668
rect 18676 17612 18686 17668
rect 16156 17556 16212 17612
rect 14466 17500 14476 17556
rect 14532 17500 16212 17556
rect 22194 17500 22204 17556
rect 22260 17500 23436 17556
rect 23492 17500 23502 17556
rect 13010 17388 13020 17444
rect 13076 17388 15148 17444
rect 15204 17388 15214 17444
rect 19506 17388 19516 17444
rect 19572 17388 21532 17444
rect 21588 17388 22316 17444
rect 22372 17388 22382 17444
rect 20738 17276 20748 17332
rect 20804 17276 22428 17332
rect 22484 17276 23100 17332
rect 23156 17276 23166 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 22530 17164 22540 17220
rect 22596 17164 23660 17220
rect 23716 17164 23726 17220
rect 20066 17052 20076 17108
rect 20132 17052 20524 17108
rect 20580 17052 21196 17108
rect 21252 17052 21262 17108
rect 21410 17052 21420 17108
rect 21476 17052 22876 17108
rect 22932 17052 22942 17108
rect 22642 16940 22652 16996
rect 22708 16940 23772 16996
rect 23828 16940 23838 16996
rect 14578 16828 14588 16884
rect 14644 16828 16716 16884
rect 16772 16828 16782 16884
rect 19282 16828 19292 16884
rect 19348 16828 22316 16884
rect 22372 16828 22382 16884
rect 22978 16828 22988 16884
rect 23044 16828 23996 16884
rect 24052 16828 24062 16884
rect 24210 16828 24220 16884
rect 24276 16828 26124 16884
rect 26180 16828 26190 16884
rect 21634 16716 21644 16772
rect 21700 16716 22428 16772
rect 22484 16716 22494 16772
rect 22754 16716 22764 16772
rect 22820 16716 23548 16772
rect 23604 16716 23614 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 18022 16268 18060 16324
rect 18116 16268 18126 16324
rect 23090 16156 23100 16212
rect 23156 16156 23996 16212
rect 24052 16156 24062 16212
rect 12450 16044 12460 16100
rect 12516 16044 15148 16100
rect 17490 16044 17500 16100
rect 17556 16044 19404 16100
rect 19460 16044 19470 16100
rect 15092 15876 15148 16044
rect 18386 15932 18396 15988
rect 18452 15932 19180 15988
rect 19236 15932 21420 15988
rect 21476 15932 21486 15988
rect 15092 15820 17276 15876
rect 17332 15820 18732 15876
rect 18788 15820 19404 15876
rect 19460 15820 19470 15876
rect 18274 15708 18284 15764
rect 18340 15708 18350 15764
rect 18284 15540 18340 15708
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 11778 15484 11788 15540
rect 11844 15484 14252 15540
rect 14308 15484 14700 15540
rect 14756 15484 15036 15540
rect 15092 15484 15102 15540
rect 18284 15484 19964 15540
rect 20020 15484 20030 15540
rect 17378 15372 17388 15428
rect 17444 15372 18732 15428
rect 18788 15372 18798 15428
rect 16594 15260 16604 15316
rect 16660 15260 17500 15316
rect 17556 15260 17566 15316
rect 18498 15260 18508 15316
rect 18564 15260 19516 15316
rect 19572 15260 20300 15316
rect 20356 15260 20366 15316
rect 21298 15260 21308 15316
rect 21364 15260 23212 15316
rect 23268 15260 24332 15316
rect 24388 15260 26460 15316
rect 26516 15260 26526 15316
rect 16706 15148 16716 15204
rect 16772 15148 18620 15204
rect 18676 15148 18686 15204
rect 24210 15148 24220 15204
rect 24276 15148 25228 15204
rect 25284 15148 25294 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 20962 14700 20972 14756
rect 21028 14700 22988 14756
rect 23044 14700 23054 14756
rect 14690 14476 14700 14532
rect 14756 14476 16380 14532
rect 16436 14476 16446 14532
rect 17938 14476 17948 14532
rect 18004 14476 18060 14532
rect 18116 14476 18126 14532
rect 19618 14252 19628 14308
rect 19684 14252 20412 14308
rect 20468 14252 20478 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 16818 13916 16828 13972
rect 16884 13916 17500 13972
rect 17556 13916 17566 13972
rect 23090 13580 23100 13636
rect 23156 13580 23884 13636
rect 23940 13580 24556 13636
rect 24612 13580 24622 13636
rect 41200 13524 42000 13552
rect 40226 13468 40236 13524
rect 40292 13468 42000 13524
rect 41200 13440 42000 13468
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 24882 5180 24892 5236
rect 24948 5180 26124 5236
rect 26180 5180 26190 5236
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 17490 4060 17500 4116
rect 17556 4060 18732 4116
rect 18788 4060 18798 4116
rect 20850 4060 20860 4116
rect 20916 4060 22092 4116
rect 22148 4060 22158 4116
rect 24210 4060 24220 4116
rect 24276 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 21522 3612 21532 3668
rect 21588 3612 22428 3668
rect 22484 3612 22494 3668
rect 23538 3612 23548 3668
rect 23604 3612 25564 3668
rect 25620 3612 25630 3668
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 19404 23436 19460 23492
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19516 20412 19572 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 19404 20076 19460 20132
rect 19516 19852 19572 19908
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 18060 16268 18116 16324
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 18060 14476 18116 14532
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 19404 23492 19460 23502
rect 19404 20132 19460 23436
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19404 20066 19460 20076
rect 19516 20468 19572 20478
rect 19516 19908 19572 20412
rect 19516 19842 19572 19852
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 18060 16324 18116 16334
rect 18060 14532 18116 16268
rect 18060 14466 18116 14476
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13888 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _102_
timestamp 1698175906
transform 1 0 15232 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15344 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform 1 0 18032 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform 1 0 14336 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform 1 0 18704 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform 1 0 17584 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20608 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 22736 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22848 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _116_
timestamp 1698175906
transform 1 0 22400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _117_
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _118_
timestamp 1698175906
transform 1 0 19712 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _119_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16912 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 16240 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 18704 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _125_
timestamp 1698175906
transform -1 0 14896 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _127_
timestamp 1698175906
transform 1 0 17920 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _128_
timestamp 1698175906
transform -1 0 14896 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _129_
timestamp 1698175906
transform 1 0 14896 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _130_
timestamp 1698175906
transform -1 0 15456 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _132_
timestamp 1698175906
transform 1 0 15568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17920 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _134_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16464 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _135_
timestamp 1698175906
transform 1 0 13664 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _136_
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _137_
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform 1 0 17360 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _139_
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform -1 0 19376 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform 1 0 19488 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _142_
timestamp 1698175906
transform -1 0 19712 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _143_
timestamp 1698175906
transform -1 0 16464 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _144_
timestamp 1698175906
transform 1 0 16576 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18480 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 21728 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _147_
timestamp 1698175906
transform 1 0 20272 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _148_
timestamp 1698175906
transform -1 0 23296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform 1 0 22064 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform -1 0 20272 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform 1 0 17808 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform -1 0 20832 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19936 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _154_
timestamp 1698175906
transform -1 0 14896 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 18816 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14672 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _158_
timestamp 1698175906
transform 1 0 13776 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14896 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_
timestamp 1698175906
transform 1 0 21392 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _161_
timestamp 1698175906
transform 1 0 15456 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _162_
timestamp 1698175906
transform 1 0 22064 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _163_
timestamp 1698175906
transform 1 0 23744 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _164_
timestamp 1698175906
transform 1 0 18480 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform 1 0 22064 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _167_
timestamp 1698175906
transform 1 0 23408 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _168_
timestamp 1698175906
transform 1 0 24192 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _169_
timestamp 1698175906
transform 1 0 25200 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform 1 0 20832 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _171_
timestamp 1698175906
transform 1 0 19488 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform 1 0 21840 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform -1 0 26544 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _174_
timestamp 1698175906
transform 1 0 25984 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _175_
timestamp 1698175906
transform 1 0 23856 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _176_
timestamp 1698175906
transform 1 0 26768 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform 1 0 21280 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _178_
timestamp 1698175906
transform 1 0 26544 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _179_
timestamp 1698175906
transform -1 0 19712 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _180_
timestamp 1698175906
transform 1 0 23296 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _181_
timestamp 1698175906
transform 1 0 18816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _182_
timestamp 1698175906
transform -1 0 23296 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _183_
timestamp 1698175906
transform 1 0 22176 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _184_
timestamp 1698175906
transform 1 0 21056 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform -1 0 17024 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 16464 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform -1 0 22736 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _188_
timestamp 1698175906
transform -1 0 20160 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform -1 0 27552 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _190_
timestamp 1698175906
transform 1 0 25760 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_
timestamp 1698175906
transform -1 0 20720 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18592 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _193_
timestamp 1698175906
transform 1 0 23856 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _194_
timestamp 1698175906
transform -1 0 25760 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _195_
timestamp 1698175906
transform -1 0 17920 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _196_
timestamp 1698175906
transform 1 0 17920 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _197_
timestamp 1698175906
transform -1 0 18368 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _198_
timestamp 1698175906
transform 1 0 18368 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _199_
timestamp 1698175906
transform -1 0 17024 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_
timestamp 1698175906
transform -1 0 27664 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _201_
timestamp 1698175906
transform 1 0 26096 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 11536 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 10416 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 9856 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 10752 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 17584 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform -1 0 15792 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 18368 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 20832 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform -1 0 14000 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 22736 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 24976 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 25648 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 23072 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 21168 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 14336 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 20160 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 17696 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform 1 0 21616 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 14448 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 25536 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _229_
timestamp 1698175906
transform 1 0 17584 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _230_
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _231_
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__A1
timestamp 1698175906
transform 1 0 14896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__A2
timestamp 1698175906
transform 1 0 27776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A2
timestamp 1698175906
transform 1 0 27888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 25984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 17472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 13664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 14224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 21392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 16016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform -1 0 21840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 24304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 14224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 27328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 23632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 25424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 26544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 18480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 24416 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 25088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform -1 0 17696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 25312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 18032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18032 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20496 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698175906
transform 1 0 17472 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_171
timestamp 1698175906
transform 1 0 20496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_201 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23856 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_209
timestamp 1698175906
transform 1 0 24752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_237
timestamp 1698175906
transform 1 0 27888 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1698175906
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_143
timestamp 1698175906
transform 1 0 17360 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_183
timestamp 1698175906
transform 1 0 21840 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_215 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25424 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698175906
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698175906
transform 1 0 28112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698175906
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_104
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_120
timestamp 1698175906
transform 1 0 14784 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_128
timestamp 1698175906
transform 1 0 15680 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_132
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_171
timestamp 1698175906
transform 1 0 20496 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_173
timestamp 1698175906
transform 1 0 20720 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_203
timestamp 1698175906
transform 1 0 24080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698175906
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_314
timestamp 1698175906
transform 1 0 36512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_330
timestamp 1698175906
transform 1 0 38304 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_338
timestamp 1698175906
transform 1 0 39200 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_342
timestamp 1698175906
transform 1 0 39648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_344
timestamp 1698175906
transform 1 0 39872 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_146
timestamp 1698175906
transform 1 0 17696 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_153
timestamp 1698175906
transform 1 0 18480 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_166
timestamp 1698175906
transform 1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_168
timestamp 1698175906
transform 1 0 20160 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_173
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_189
timestamp 1698175906
transform 1 0 22512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_191
timestamp 1698175906
transform 1 0 22736 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_196
timestamp 1698175906
transform 1 0 23296 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_228
timestamp 1698175906
transform 1 0 26880 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_88
timestamp 1698175906
transform 1 0 11200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_90
timestamp 1698175906
transform 1 0 11424 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_124
timestamp 1698175906
transform 1 0 15232 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_160
timestamp 1698175906
transform 1 0 19264 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_164
timestamp 1698175906
transform 1 0 19712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_139
timestamp 1698175906
transform 1 0 16912 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_154
timestamp 1698175906
transform 1 0 18592 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_164
timestamp 1698175906
transform 1 0 19712 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_193
timestamp 1698175906
transform 1 0 22960 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_223
timestamp 1698175906
transform 1 0 26320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_227
timestamp 1698175906
transform 1 0 26768 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 10304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_113
timestamp 1698175906
transform 1 0 14000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_117
timestamp 1698175906
transform 1 0 14448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698175906
transform 1 0 16240 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_174
timestamp 1698175906
transform 1 0 20832 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_109
timestamp 1698175906
transform 1 0 13552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_112
timestamp 1698175906
transform 1 0 13888 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_114
timestamp 1698175906
transform 1 0 14112 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_145
timestamp 1698175906
transform 1 0 17584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_149
timestamp 1698175906
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_151
timestamp 1698175906
transform 1 0 18256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698175906
transform 1 0 20384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_185
timestamp 1698175906
transform 1 0 22064 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_196
timestamp 1698175906
transform 1 0 23296 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_228
timestamp 1698175906
transform 1 0 26880 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 4480 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_80
timestamp 1698175906
transform 1 0 10304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_110
timestamp 1698175906
transform 1 0 13664 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_158
timestamp 1698175906
transform 1 0 19040 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_179
timestamp 1698175906
transform 1 0 21392 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_195
timestamp 1698175906
transform 1 0 23184 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698175906
transform 1 0 24080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_207
timestamp 1698175906
transform 1 0 24528 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_241
timestamp 1698175906
transform 1 0 28336 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698175906
transform 1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 40320 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_191
timestamp 1698175906
transform 1 0 22736 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1698175906
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_108
timestamp 1698175906
transform 1 0 13440 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_114
timestamp 1698175906
transform 1 0 14112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_135
timestamp 1698175906
transform 1 0 16464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_148
timestamp 1698175906
transform 1 0 17920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_174
timestamp 1698175906
transform 1 0 20832 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_188
timestamp 1698175906
transform 1 0 22400 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_227
timestamp 1698175906
transform 1 0 26768 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_259
timestamp 1698175906
transform 1 0 30352 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698175906
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_119
timestamp 1698175906
transform 1 0 14672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698175906
transform 1 0 15120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_125
timestamp 1698175906
transform 1 0 15344 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_139
timestamp 1698175906
transform 1 0 16912 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_161
timestamp 1698175906
transform 1 0 19376 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_230
timestamp 1698175906
transform 1 0 27104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_234
timestamp 1698175906
transform 1 0 27552 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_113
timestamp 1698175906
transform 1 0 14000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_117
timestamp 1698175906
transform 1 0 14448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_135
timestamp 1698175906
transform 1 0 16464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_199
timestamp 1698175906
transform 1 0 23632 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_214
timestamp 1698175906
transform 1 0 25312 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_246
timestamp 1698175906
transform 1 0 28896 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 9072 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698175906
transform 1 0 9744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_111
timestamp 1698175906
transform 1 0 13776 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_122
timestamp 1698175906
transform 1 0 15008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_124
timestamp 1698175906
transform 1 0 15232 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_148
timestamp 1698175906
transform 1 0 17920 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_152
timestamp 1698175906
transform 1 0 18368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_154
timestamp 1698175906
transform 1 0 18592 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_161
timestamp 1698175906
transform 1 0 19376 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_169
timestamp 1698175906
transform 1 0 20272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698175906
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_234
timestamp 1698175906
transform 1 0 27552 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698175906
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_120
timestamp 1698175906
transform 1 0 14784 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_128
timestamp 1698175906
transform 1 0 15680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698175906
transform 1 0 17472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_151
timestamp 1698175906
transform 1 0 18256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_204
timestamp 1698175906
transform 1 0 24192 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698175906
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_220
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_229
timestamp 1698175906
transform 1 0 26992 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_235
timestamp 1698175906
transform 1 0 27664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_239
timestamp 1698175906
transform 1 0 28112 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_271
timestamp 1698175906
transform 1 0 31696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_131
timestamp 1698175906
transform 1 0 16016 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698175906
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_142
timestamp 1698175906
transform 1 0 17248 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_149
timestamp 1698175906
transform 1 0 18032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_159
timestamp 1698175906
transform 1 0 19152 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_185
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_197
timestamp 1698175906
transform 1 0 23408 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_213
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_104
timestamp 1698175906
transform 1 0 12992 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_112
timestamp 1698175906
transform 1 0 13888 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_116
timestamp 1698175906
transform 1 0 14336 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_121
timestamp 1698175906
transform 1 0 14896 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_155
timestamp 1698175906
transform 1 0 18704 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_171
timestamp 1698175906
transform 1 0 20496 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_180
timestamp 1698175906
transform 1 0 21504 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_184
timestamp 1698175906
transform 1 0 21952 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_190
timestamp 1698175906
transform 1 0 22624 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_142
timestamp 1698175906
transform 1 0 17248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_146
timestamp 1698175906
transform 1 0 17696 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_162
timestamp 1698175906
transform 1 0 19488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_170
timestamp 1698175906
transform 1 0 20384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_209
timestamp 1698175906
transform 1 0 24752 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_211
timestamp 1698175906
transform 1 0 24976 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_214
timestamp 1698175906
transform 1 0 25312 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_226
timestamp 1698175906
transform 1 0 26656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_228
timestamp 1698175906
transform 1 0 26880 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_234
timestamp 1698175906
transform 1 0 27552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_96
timestamp 1698175906
transform 1 0 12096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_129
timestamp 1698175906
transform 1 0 15792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698175906
transform 1 0 16240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_137
timestamp 1698175906
transform 1 0 16688 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_148
timestamp 1698175906
transform 1 0 17920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_152
timestamp 1698175906
transform 1 0 18368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_154
timestamp 1698175906
transform 1 0 18592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_177
timestamp 1698175906
transform 1 0 21168 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_181
timestamp 1698175906
transform 1 0 21616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_185
timestamp 1698175906
transform 1 0 22064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_187
timestamp 1698175906
transform 1 0 22288 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_243
timestamp 1698175906
transform 1 0 28560 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_275
timestamp 1698175906
transform 1 0 32144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_139
timestamp 1698175906
transform 1 0 16912 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_143
timestamp 1698175906
transform 1 0 17360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_182
timestamp 1698175906
transform 1 0 21728 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_184
timestamp 1698175906
transform 1 0 21952 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_218
timestamp 1698175906
transform 1 0 25760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_222
timestamp 1698175906
transform 1 0 26208 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_128
timestamp 1698175906
transform 1 0 15680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_148
timestamp 1698175906
transform 1 0 17920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_216
timestamp 1698175906
transform 1 0 25536 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_115
timestamp 1698175906
transform 1 0 14224 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_151
timestamp 1698175906
transform 1 0 18256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_155
timestamp 1698175906
transform 1 0 18704 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_183
timestamp 1698175906
transform 1 0 21840 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_215
timestamp 1698175906
transform 1 0 25424 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_231
timestamp 1698175906
transform 1 0 27216 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_239
timestamp 1698175906
transform 1 0 28112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698175906
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698175906
transform 1 0 19824 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 24080 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698175906
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698175906
transform 1 0 23856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_203
timestamp 1698175906
transform 1 0 24080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita56_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 27776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita56_26
timestamp 1698175906
transform 1 0 39984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20944 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 24976 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 16912 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 17584 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 4480 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 21280 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 17360 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 20272 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform -1 0 4480 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 26208 41200 26320 42000 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 41200 13440 42000 13552 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 20160 41200 20272 42000 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 24192 42000 24304 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 24192 41200 24304 42000 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 26040 19488 26040 19488 0 _000_
rlabel metal2 24808 19208 24808 19208 0 _001_
rlabel metal2 26824 21224 26824 21224 0 _002_
rlabel metal3 23576 16184 23576 16184 0 _003_
rlabel metal2 22064 15400 22064 15400 0 _004_
rlabel metal2 15960 28280 15960 28280 0 _005_
rlabel metal3 20496 23128 20496 23128 0 _006_
rlabel metal2 26040 25872 26040 25872 0 _007_
rlabel metal2 18648 13272 18648 13272 0 _008_
rlabel metal2 25480 27496 25480 27496 0 _009_
rlabel metal2 18144 13832 18144 13832 0 _010_
rlabel metal2 15400 14840 15400 14840 0 _011_
rlabel metal2 26432 23352 26432 23352 0 _012_
rlabel metal2 22848 26936 22848 26936 0 _013_
rlabel metal2 14616 25144 14616 25144 0 _014_
rlabel metal2 12488 15736 12488 15736 0 _015_
rlabel metal3 12656 18312 12656 18312 0 _016_
rlabel metal2 10808 21952 10808 21952 0 _017_
rlabel metal2 11704 21784 11704 21784 0 _018_
rlabel metal2 18704 26936 18704 26936 0 _019_
rlabel metal2 14840 25928 14840 25928 0 _020_
rlabel metal2 20552 26656 20552 26656 0 _021_
rlabel metal2 21448 15512 21448 15512 0 _022_
rlabel metal2 13048 17192 13048 17192 0 _023_
rlabel metal2 23688 21896 23688 21896 0 _024_
rlabel metal2 18088 17640 18088 17640 0 _025_
rlabel metal2 19488 14392 19488 14392 0 _026_
rlabel metal3 20888 17080 20888 17080 0 _027_
rlabel metal2 14616 18312 14616 18312 0 _028_
rlabel metal2 18816 14728 18816 14728 0 _029_
rlabel metal2 15064 17976 15064 17976 0 _030_
rlabel metal2 16464 18312 16464 18312 0 _031_
rlabel metal2 14504 17976 14504 17976 0 _032_
rlabel metal2 27160 21168 27160 21168 0 _033_
rlabel metal2 22232 20832 22232 20832 0 _034_
rlabel metal3 20832 16856 20832 16856 0 _035_
rlabel metal2 24024 22344 24024 22344 0 _036_
rlabel metal2 22232 24640 22232 24640 0 _037_
rlabel metal3 24248 24920 24248 24920 0 _038_
rlabel metal2 23576 23296 23576 23296 0 _039_
rlabel metal2 26824 22400 26824 22400 0 _040_
rlabel metal2 25928 20496 25928 20496 0 _041_
rlabel metal2 21448 19712 21448 19712 0 _042_
rlabel metal3 21112 20104 21112 20104 0 _043_
rlabel metal2 22344 20384 22344 20384 0 _044_
rlabel metal2 24584 19432 24584 19432 0 _045_
rlabel metal2 26936 21336 26936 21336 0 _046_
rlabel metal2 21784 20216 21784 20216 0 _047_
rlabel metal2 19040 14728 19040 14728 0 _048_
rlabel metal2 22792 17136 22792 17136 0 _049_
rlabel metal2 21560 17192 21560 17192 0 _050_
rlabel metal2 21672 16856 21672 16856 0 _051_
rlabel metal2 16408 27832 16408 27832 0 _052_
rlabel metal2 20104 23240 20104 23240 0 _053_
rlabel metal2 26824 25480 26824 25480 0 _054_
rlabel metal3 20048 14280 20048 14280 0 _055_
rlabel metal3 24976 26936 24976 26936 0 _056_
rlabel metal2 17584 15064 17584 15064 0 _057_
rlabel metal2 17696 15288 17696 15288 0 _058_
rlabel metal3 17696 15176 17696 15176 0 _059_
rlabel metal2 27048 23128 27048 23128 0 _060_
rlabel metal2 15064 21952 15064 21952 0 _061_
rlabel metal2 15512 22624 15512 22624 0 _062_
rlabel metal2 27384 25760 27384 25760 0 _063_
rlabel metal3 22568 26936 22568 26936 0 _064_
rlabel metal2 13832 18592 13832 18592 0 _065_
rlabel metal2 21224 24752 21224 24752 0 _066_
rlabel metal2 14840 21056 14840 21056 0 _067_
rlabel metal2 19208 21448 19208 21448 0 _068_
rlabel metal2 17640 23856 17640 23856 0 _069_
rlabel metal2 18088 23520 18088 23520 0 _070_
rlabel metal2 21336 25536 21336 25536 0 _071_
rlabel metal3 19432 18424 19432 18424 0 _072_
rlabel metal2 21672 20104 21672 20104 0 _073_
rlabel metal2 26152 25088 26152 25088 0 _074_
rlabel metal2 22680 26264 22680 26264 0 _075_
rlabel metal3 18200 20104 18200 20104 0 _076_
rlabel metal2 21560 21168 21560 21168 0 _077_
rlabel metal3 16184 20104 16184 20104 0 _078_
rlabel metal3 18592 21336 18592 21336 0 _079_
rlabel metal2 16968 23800 16968 23800 0 _080_
rlabel metal2 18872 24248 18872 24248 0 _081_
rlabel metal2 16632 24360 16632 24360 0 _082_
rlabel metal2 14728 24360 14728 24360 0 _083_
rlabel metal2 14728 18088 14728 18088 0 _084_
rlabel metal2 18536 19992 18536 19992 0 _085_
rlabel metal2 14728 19264 14728 19264 0 _086_
rlabel metal2 16128 27944 16128 27944 0 _087_
rlabel metal2 16520 20888 16520 20888 0 _088_
rlabel metal2 13944 19600 13944 19600 0 _089_
rlabel metal3 18480 16072 18480 16072 0 _090_
rlabel metal2 21392 19208 21392 19208 0 _091_
rlabel metal3 18760 24920 18760 24920 0 _092_
rlabel metal2 19432 26040 19432 26040 0 _093_
rlabel metal2 20104 18648 20104 18648 0 _094_
rlabel metal2 17136 25480 17136 25480 0 _095_
rlabel metal2 16184 25144 16184 25144 0 _096_
rlabel metal2 19656 23688 19656 23688 0 _097_
rlabel metal2 21224 26544 21224 26544 0 _098_
rlabel metal3 22008 14728 22008 14728 0 _099_
rlabel metal2 23128 17360 23128 17360 0 _100_
rlabel metal3 2478 28280 2478 28280 0 clk
rlabel metal2 20328 20888 20328 20888 0 clknet_0_clk
rlabel metal3 18032 28616 18032 28616 0 clknet_1_0__leaf_clk
rlabel metal2 21784 28224 21784 28224 0 clknet_1_1__leaf_clk
rlabel metal2 14616 16016 14616 16016 0 dut56.count\[0\]
rlabel metal2 13496 19264 13496 19264 0 dut56.count\[1\]
rlabel metal3 13496 22456 13496 22456 0 dut56.count\[2\]
rlabel metal2 13832 20804 13832 20804 0 dut56.count\[3\]
rlabel metal2 21112 6356 21112 6356 0 net1
rlabel metal2 17752 6356 17752 6356 0 net10
rlabel metal2 37912 21672 37912 21672 0 net11
rlabel metal2 28168 18704 28168 18704 0 net12
rlabel metal2 4312 18032 4312 18032 0 net13
rlabel metal2 27272 25760 27272 25760 0 net14
rlabel metal2 21448 5964 21448 5964 0 net15
rlabel metal3 24248 13608 24248 13608 0 net16
rlabel metal2 21448 27328 21448 27328 0 net17
rlabel metal2 17696 28056 17696 28056 0 net18
rlabel metal2 12712 26208 12712 26208 0 net19
rlabel metal3 29988 19320 29988 19320 0 net2
rlabel metal2 20664 32200 20664 32200 0 net20
rlabel metal3 31920 23184 31920 23184 0 net21
rlabel metal2 4312 25424 4312 25424 0 net22
rlabel metal2 27384 23688 27384 23688 0 net23
rlabel metal2 25088 38024 25088 38024 0 net24
rlabel metal3 26880 37912 26880 37912 0 net25
rlabel metal2 40264 13664 40264 13664 0 net26
rlabel metal2 25368 6748 25368 6748 0 net3
rlabel metal2 24192 15176 24192 15176 0 net4
rlabel metal2 27384 21784 27384 21784 0 net5
rlabel metal2 18088 30212 18088 30212 0 net6
rlabel metal2 24696 28112 24696 28112 0 net7
rlabel metal2 17416 28392 17416 28392 0 net8
rlabel metal2 20216 13944 20216 13944 0 net9
rlabel metal2 20888 2422 20888 2422 0 segm[0]
rlabel metal2 40040 19656 40040 19656 0 segm[10]
rlabel metal2 24920 2982 24920 2982 0 segm[11]
rlabel metal2 24248 2422 24248 2422 0 segm[12]
rlabel metal2 40040 21504 40040 21504 0 segm[13]
rlabel metal2 18200 39746 18200 39746 0 segm[1]
rlabel metal2 24920 39354 24920 39354 0 segm[3]
rlabel metal2 16856 38962 16856 38962 0 segm[4]
rlabel metal2 18200 2198 18200 2198 0 segm[6]
rlabel metal2 17528 2422 17528 2422 0 segm[7]
rlabel metal2 40040 22344 40040 22344 0 segm[8]
rlabel metal2 40040 19096 40040 19096 0 segm[9]
rlabel metal3 1358 18200 1358 18200 0 sel[0]
rlabel metal2 40040 26712 40040 26712 0 sel[10]
rlabel metal2 21560 2198 21560 2198 0 sel[11]
rlabel metal2 23576 2198 23576 2198 0 sel[1]
rlabel metal2 20888 39746 20888 39746 0 sel[2]
rlabel metal2 17528 39354 17528 39354 0 sel[3]
rlabel metal3 1358 25592 1358 25592 0 sel[4]
rlabel metal2 20216 39354 20216 39354 0 sel[5]
rlabel metal3 40642 22904 40642 22904 0 sel[6]
rlabel metal3 1414 24920 1414 24920 0 sel[7]
rlabel metal2 40040 24360 40040 24360 0 sel[8]
rlabel metal2 24248 39746 24248 39746 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
