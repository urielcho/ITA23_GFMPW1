magic
tech gf180mcuD
magscale 1 5
timestamp 1699641800
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 9408 20600 9464 21000
rect 10416 20600 10472 21000
rect 11088 20600 11144 21000
rect 12432 20600 12488 21000
rect 8400 0 8456 400
<< obsm2 >>
rect 966 20570 9378 20600
rect 9494 20570 10386 20600
rect 10502 20570 11058 20600
rect 11174 20570 12402 20600
rect 12518 20570 20146 20600
rect 966 430 20146 20570
rect 966 400 8370 430
rect 8486 400 20146 430
<< metal3 >>
rect 20600 18480 21000 18536
rect 20600 13440 21000 13496
rect 0 13104 400 13160
rect 20600 13104 21000 13160
rect 0 12768 400 12824
rect 20600 12768 21000 12824
rect 0 12432 400 12488
rect 20600 12432 21000 12488
rect 0 12096 400 12152
rect 20600 12096 21000 12152
rect 20600 11760 21000 11816
rect 20600 11424 21000 11480
rect 20600 11088 21000 11144
rect 0 10752 400 10808
rect 20600 10752 21000 10808
rect 0 9744 400 9800
rect 20600 9744 21000 9800
rect 20600 9408 21000 9464
rect 20600 9072 21000 9128
rect 0 8736 400 8792
rect 20600 8736 21000 8792
rect 0 8400 400 8456
<< obsm3 >>
rect 400 18566 20600 19222
rect 400 18450 20570 18566
rect 400 13526 20600 18450
rect 400 13410 20570 13526
rect 400 13190 20600 13410
rect 430 13074 20570 13190
rect 400 12854 20600 13074
rect 430 12738 20570 12854
rect 400 12518 20600 12738
rect 430 12402 20570 12518
rect 400 12182 20600 12402
rect 430 12066 20570 12182
rect 400 11846 20600 12066
rect 400 11730 20570 11846
rect 400 11510 20600 11730
rect 400 11394 20570 11510
rect 400 11174 20600 11394
rect 400 11058 20570 11174
rect 400 10838 20600 11058
rect 430 10722 20570 10838
rect 400 9830 20600 10722
rect 430 9714 20570 9830
rect 400 9494 20600 9714
rect 400 9378 20570 9494
rect 400 9158 20600 9378
rect 400 9042 20570 9158
rect 400 8822 20600 9042
rect 430 8706 20570 8822
rect 400 8486 20600 8706
rect 430 8370 20600 8486
rect 400 1554 20600 8370
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 10654 8913 10682 9791
<< labels >>
rlabel metal3 s 0 12096 400 12152 6 clk
port 1 nsew signal input
rlabel metal3 s 20600 18480 21000 18536 6 segm[0]
port 2 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 segm[10]
port 3 nsew signal output
rlabel metal3 s 20600 11088 21000 11144 6 segm[11]
port 4 nsew signal output
rlabel metal3 s 20600 10752 21000 10808 6 segm[12]
port 5 nsew signal output
rlabel metal2 s 9408 20600 9464 21000 6 segm[13]
port 6 nsew signal output
rlabel metal3 s 0 13104 400 13160 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 20600 13440 21000 13496 6 segm[2]
port 8 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 segm[3]
port 9 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 segm[4]
port 10 nsew signal output
rlabel metal2 s 10416 20600 10472 21000 6 segm[5]
port 11 nsew signal output
rlabel metal3 s 20600 12096 21000 12152 6 segm[6]
port 12 nsew signal output
rlabel metal3 s 20600 9408 21000 9464 6 segm[7]
port 13 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 20600 9744 21000 9800 6 segm[9]
port 15 nsew signal output
rlabel metal2 s 11088 20600 11144 21000 6 sel[0]
port 16 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 sel[10]
port 17 nsew signal output
rlabel metal3 s 0 10752 400 10808 6 sel[11]
port 18 nsew signal output
rlabel metal2 s 12432 20600 12488 21000 6 sel[1]
port 19 nsew signal output
rlabel metal3 s 20600 11760 21000 11816 6 sel[2]
port 20 nsew signal output
rlabel metal3 s 20600 13104 21000 13160 6 sel[3]
port 21 nsew signal output
rlabel metal3 s 20600 12768 21000 12824 6 sel[4]
port 22 nsew signal output
rlabel metal3 s 0 12432 400 12488 6 sel[5]
port 23 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 sel[6]
port 24 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 sel[7]
port 25 nsew signal output
rlabel metal3 s 20600 11424 21000 11480 6 sel[8]
port 26 nsew signal output
rlabel metal3 s 20600 8736 21000 8792 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 459948
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita54/runs/23_11_10_12_41/results/signoff/ita54.magic.gds
string GDS_START 150106
<< end >>

