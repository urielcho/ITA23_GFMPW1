magic
tech gf180mcuD
magscale 1 5
timestamp 1699645780
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 8801 18999 8807 19025
rect 8833 18999 8839 19025
rect 10705 18999 10711 19025
rect 10737 18999 10743 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 3151 18969 3177 18975
rect 3151 18937 3177 18943
rect 10487 18969 10513 18975
rect 10487 18937 10513 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9199 18745 9225 18751
rect 9199 18713 9225 18719
rect 10711 18745 10737 18751
rect 10711 18713 10737 18719
rect 8689 18607 8695 18633
rect 8721 18607 8727 18633
rect 10201 18607 10207 18633
rect 10233 18607 10239 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 9927 14265 9953 14271
rect 9927 14233 9953 14239
rect 9983 14265 10009 14271
rect 9983 14233 10009 14239
rect 10263 14265 10289 14271
rect 10263 14233 10289 14239
rect 10319 14265 10345 14271
rect 10319 14233 10345 14239
rect 9815 14209 9841 14215
rect 9815 14177 9841 14183
rect 10431 14209 10457 14215
rect 10431 14177 10457 14183
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8751 14041 8777 14047
rect 8751 14009 8777 14015
rect 8807 13985 8833 13991
rect 8807 13953 8833 13959
rect 8639 13929 8665 13935
rect 7009 13903 7015 13929
rect 7041 13903 7047 13929
rect 9585 13903 9591 13929
rect 9617 13903 9623 13929
rect 8639 13897 8665 13903
rect 9087 13873 9113 13879
rect 7345 13847 7351 13873
rect 7377 13847 7383 13873
rect 8409 13847 8415 13873
rect 8441 13847 8447 13873
rect 9087 13841 9113 13847
rect 9479 13873 9505 13879
rect 9977 13847 9983 13873
rect 10009 13847 10015 13873
rect 11041 13847 11047 13873
rect 11073 13847 11079 13873
rect 9479 13841 9505 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 8527 13593 8553 13599
rect 20007 13593 20033 13599
rect 8185 13567 8191 13593
rect 8217 13567 8223 13593
rect 10369 13567 10375 13593
rect 10401 13567 10407 13593
rect 10817 13567 10823 13593
rect 10849 13567 10855 13593
rect 8527 13561 8553 13567
rect 20007 13561 20033 13567
rect 8639 13537 8665 13543
rect 6785 13511 6791 13537
rect 6817 13511 6823 13537
rect 8913 13511 8919 13537
rect 8945 13511 8951 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 8639 13505 8665 13511
rect 8471 13481 8497 13487
rect 7121 13455 7127 13481
rect 7153 13455 7159 13481
rect 8471 13449 8497 13455
rect 8751 13481 8777 13487
rect 10655 13481 10681 13487
rect 9305 13455 9311 13481
rect 9337 13455 9343 13481
rect 8751 13449 8777 13455
rect 10655 13449 10681 13455
rect 10767 13425 10793 13431
rect 10767 13393 10793 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7631 13257 7657 13263
rect 7631 13225 7657 13231
rect 8751 13257 8777 13263
rect 8751 13225 8777 13231
rect 9591 13257 9617 13263
rect 9591 13225 9617 13231
rect 10039 13257 10065 13263
rect 10039 13225 10065 13231
rect 8023 13201 8049 13207
rect 8023 13169 8049 13175
rect 8191 13201 8217 13207
rect 8191 13169 8217 13175
rect 8975 13201 9001 13207
rect 8975 13169 9001 13175
rect 9703 13201 9729 13207
rect 9703 13169 9729 13175
rect 9815 13201 9841 13207
rect 9815 13169 9841 13175
rect 10151 13201 10177 13207
rect 10151 13169 10177 13175
rect 10263 13201 10289 13207
rect 13063 13201 13089 13207
rect 10873 13175 10879 13201
rect 10905 13175 10911 13201
rect 10263 13169 10289 13175
rect 13063 13169 13089 13175
rect 8303 13145 8329 13151
rect 9535 13145 9561 13151
rect 7513 13119 7519 13145
rect 7545 13119 7551 13145
rect 9081 13119 9087 13145
rect 9113 13119 9119 13145
rect 8303 13113 8329 13119
rect 9535 13113 9561 13119
rect 9927 13145 9953 13151
rect 10537 13119 10543 13145
rect 10569 13119 10575 13145
rect 12833 13119 12839 13145
rect 12865 13119 12871 13145
rect 12945 13119 12951 13145
rect 12977 13119 12983 13145
rect 18937 13119 18943 13145
rect 18969 13119 18975 13145
rect 9927 13113 9953 13119
rect 8079 13089 8105 13095
rect 12223 13089 12249 13095
rect 11937 13063 11943 13089
rect 11969 13063 11975 13089
rect 8079 13057 8105 13063
rect 12223 13057 12249 13063
rect 13679 13089 13705 13095
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 13679 13057 13705 13063
rect 7687 13033 7713 13039
rect 7687 13001 7713 13007
rect 12895 13033 12921 13039
rect 12895 13001 12921 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 967 12809 993 12815
rect 967 12777 993 12783
rect 8303 12809 8329 12815
rect 20007 12809 20033 12815
rect 10761 12783 10767 12809
rect 10793 12783 10799 12809
rect 13505 12783 13511 12809
rect 13537 12783 13543 12809
rect 8303 12777 8329 12783
rect 20007 12777 20033 12783
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 10985 12727 10991 12753
rect 11017 12727 11023 12753
rect 12105 12727 12111 12753
rect 12137 12727 12143 12753
rect 14177 12727 14183 12753
rect 14209 12727 14215 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 13791 12697 13817 12703
rect 8521 12671 8527 12697
rect 8553 12671 8559 12697
rect 12441 12671 12447 12697
rect 12473 12671 12479 12697
rect 14289 12671 14295 12697
rect 14321 12671 14327 12697
rect 13791 12665 13817 12671
rect 8695 12641 8721 12647
rect 8695 12609 8721 12615
rect 10711 12641 10737 12647
rect 10711 12609 10737 12615
rect 10767 12641 10793 12647
rect 10767 12609 10793 12615
rect 10879 12641 10905 12647
rect 10879 12609 10905 12615
rect 13623 12641 13649 12647
rect 13623 12609 13649 12615
rect 13735 12641 13761 12647
rect 13735 12609 13761 12615
rect 14575 12641 14601 12647
rect 14737 12615 14743 12641
rect 14769 12615 14775 12641
rect 14575 12609 14601 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 8191 12473 8217 12479
rect 8191 12441 8217 12447
rect 9871 12473 9897 12479
rect 9871 12441 9897 12447
rect 12783 12473 12809 12479
rect 12783 12441 12809 12447
rect 8919 12417 8945 12423
rect 8919 12385 8945 12391
rect 9927 12417 9953 12423
rect 13393 12391 13399 12417
rect 13425 12391 13431 12417
rect 9927 12385 9953 12391
rect 7961 12335 7967 12361
rect 7993 12335 7999 12361
rect 8689 12335 8695 12361
rect 8721 12335 8727 12361
rect 8801 12335 8807 12361
rect 8833 12335 8839 12361
rect 10033 12335 10039 12361
rect 10065 12335 10071 12361
rect 10145 12335 10151 12361
rect 10177 12335 10183 12361
rect 13001 12335 13007 12361
rect 13033 12335 13039 12361
rect 18825 12335 18831 12361
rect 18857 12335 18863 12361
rect 8751 12305 8777 12311
rect 14799 12305 14825 12311
rect 6505 12279 6511 12305
rect 6537 12279 6543 12305
rect 7569 12279 7575 12305
rect 7601 12279 7607 12305
rect 14513 12279 14519 12305
rect 14545 12279 14551 12305
rect 8751 12273 8777 12279
rect 14799 12273 14825 12279
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 7575 12081 7601 12087
rect 7575 12049 7601 12055
rect 20007 12025 20033 12031
rect 8185 11999 8191 12025
rect 8217 11999 8223 12025
rect 9529 11999 9535 12025
rect 9561 11999 9567 12025
rect 12665 11999 12671 12025
rect 12697 11999 12703 12025
rect 13337 11999 13343 12025
rect 13369 11999 13375 12025
rect 20007 11993 20033 11999
rect 7743 11969 7769 11975
rect 8247 11969 8273 11975
rect 8129 11943 8135 11969
rect 8161 11943 8167 11969
rect 7743 11937 7769 11943
rect 8247 11937 8273 11943
rect 8359 11969 8385 11975
rect 10095 11969 10121 11975
rect 12783 11969 12809 11975
rect 8465 11943 8471 11969
rect 8497 11943 8503 11969
rect 11265 11943 11271 11969
rect 11297 11943 11303 11969
rect 8359 11937 8385 11943
rect 10095 11937 10121 11943
rect 12783 11937 12809 11943
rect 12951 11969 12977 11975
rect 13169 11943 13175 11969
rect 13201 11943 13207 11969
rect 13281 11943 13287 11969
rect 13313 11943 13319 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 12951 11937 12977 11943
rect 7631 11913 7657 11919
rect 9535 11913 9561 11919
rect 9473 11887 9479 11913
rect 9505 11887 9511 11913
rect 7631 11881 7657 11887
rect 9535 11881 9561 11887
rect 9591 11913 9617 11919
rect 13399 11913 13425 11919
rect 11601 11887 11607 11913
rect 11633 11887 11639 11913
rect 9591 11881 9617 11887
rect 13399 11881 13425 11887
rect 9703 11857 9729 11863
rect 9703 11825 9729 11831
rect 10151 11857 10177 11863
rect 10151 11825 10177 11831
rect 10263 11857 10289 11863
rect 10263 11825 10289 11831
rect 12895 11857 12921 11863
rect 12895 11825 12921 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 8023 11689 8049 11695
rect 11775 11689 11801 11695
rect 9361 11663 9367 11689
rect 9393 11663 9399 11689
rect 10537 11663 10543 11689
rect 10569 11663 10575 11689
rect 8023 11657 8049 11663
rect 11775 11657 11801 11663
rect 12671 11689 12697 11695
rect 12671 11657 12697 11663
rect 12951 11689 12977 11695
rect 12951 11657 12977 11663
rect 7575 11633 7601 11639
rect 7575 11601 7601 11607
rect 9143 11633 9169 11639
rect 9143 11601 9169 11607
rect 9199 11633 9225 11639
rect 9199 11601 9225 11607
rect 10095 11633 10121 11639
rect 12727 11633 12753 11639
rect 10369 11607 10375 11633
rect 10401 11607 10407 11633
rect 10649 11607 10655 11633
rect 10681 11607 10687 11633
rect 10095 11601 10121 11607
rect 12727 11601 12753 11607
rect 7743 11577 7769 11583
rect 8247 11577 8273 11583
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 7345 11551 7351 11577
rect 7377 11551 7383 11577
rect 7905 11551 7911 11577
rect 7937 11551 7943 11577
rect 7743 11545 7769 11551
rect 8247 11545 8273 11551
rect 9031 11577 9057 11583
rect 9031 11545 9057 11551
rect 9535 11577 9561 11583
rect 9535 11545 9561 11551
rect 9703 11577 9729 11583
rect 9703 11545 9729 11551
rect 9927 11577 9953 11583
rect 11551 11577 11577 11583
rect 10817 11551 10823 11577
rect 10849 11551 10855 11577
rect 9927 11545 9953 11551
rect 11551 11545 11577 11551
rect 11719 11577 11745 11583
rect 11719 11545 11745 11551
rect 11887 11577 11913 11583
rect 11887 11545 11913 11551
rect 12559 11577 12585 11583
rect 12559 11545 12585 11551
rect 8135 11521 8161 11527
rect 5889 11495 5895 11521
rect 5921 11495 5927 11521
rect 6953 11495 6959 11521
rect 6985 11495 6991 11521
rect 8135 11489 8161 11495
rect 967 11465 993 11471
rect 967 11433 993 11439
rect 8023 11465 8049 11471
rect 8023 11433 8049 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 7407 11297 7433 11303
rect 7407 11265 7433 11271
rect 7575 11297 7601 11303
rect 7575 11265 7601 11271
rect 7967 11297 7993 11303
rect 7967 11265 7993 11271
rect 13063 11297 13089 11303
rect 13063 11265 13089 11271
rect 20007 11241 20033 11247
rect 11377 11215 11383 11241
rect 11409 11215 11415 11241
rect 20007 11209 20033 11215
rect 9479 11185 9505 11191
rect 13119 11185 13145 11191
rect 9585 11159 9591 11185
rect 9617 11159 9623 11185
rect 10649 11159 10655 11185
rect 10681 11159 10687 11185
rect 12833 11159 12839 11185
rect 12865 11159 12871 11185
rect 9479 11153 9505 11159
rect 13119 11153 13145 11159
rect 13231 11185 13257 11191
rect 13231 11153 13257 11159
rect 13287 11185 13313 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13287 11153 13313 11159
rect 7911 11129 7937 11135
rect 7911 11097 7937 11103
rect 9871 11129 9897 11135
rect 13007 11129 13033 11135
rect 10761 11103 10767 11129
rect 10793 11103 10799 11129
rect 11097 11103 11103 11129
rect 11129 11103 11135 11129
rect 12441 11103 12447 11129
rect 12473 11103 12479 11129
rect 9871 11097 9897 11103
rect 13007 11097 13033 11103
rect 7463 11073 7489 11079
rect 7463 11041 7489 11047
rect 7967 11073 7993 11079
rect 14295 11073 14321 11079
rect 9361 11047 9367 11073
rect 9393 11047 9399 11073
rect 10929 11047 10935 11073
rect 10961 11047 10967 11073
rect 7967 11041 7993 11047
rect 14295 11041 14321 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 9809 10879 9815 10905
rect 9841 10879 9847 10905
rect 8415 10849 8441 10855
rect 8415 10817 8441 10823
rect 9143 10849 9169 10855
rect 11999 10849 12025 10855
rect 9753 10823 9759 10849
rect 9785 10823 9791 10849
rect 11601 10823 11607 10849
rect 11633 10823 11639 10849
rect 13225 10823 13231 10849
rect 13257 10823 13263 10849
rect 9143 10817 9169 10823
rect 11999 10817 12025 10823
rect 7799 10793 7825 10799
rect 11775 10793 11801 10799
rect 7177 10767 7183 10793
rect 7209 10767 7215 10793
rect 8185 10767 8191 10793
rect 8217 10767 8223 10793
rect 8297 10767 8303 10793
rect 8329 10767 8335 10793
rect 8913 10767 8919 10793
rect 8945 10767 8951 10793
rect 9809 10767 9815 10793
rect 9841 10767 9847 10793
rect 10481 10767 10487 10793
rect 10513 10767 10519 10793
rect 11153 10767 11159 10793
rect 11185 10767 11191 10793
rect 7799 10761 7825 10767
rect 11775 10761 11801 10767
rect 12055 10793 12081 10799
rect 12833 10767 12839 10793
rect 12865 10767 12871 10793
rect 14513 10767 14519 10793
rect 14545 10767 14551 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 12055 10761 12081 10767
rect 6847 10737 6873 10743
rect 7289 10711 7295 10737
rect 7321 10711 7327 10737
rect 7569 10711 7575 10737
rect 7601 10711 7607 10737
rect 8353 10711 8359 10737
rect 8385 10711 8391 10737
rect 14289 10711 14295 10737
rect 14321 10711 14327 10737
rect 14849 10711 14855 10737
rect 14881 10711 14887 10737
rect 15913 10711 15919 10737
rect 15945 10711 15951 10737
rect 6847 10705 6873 10711
rect 11999 10681 12025 10687
rect 11999 10649 12025 10655
rect 20007 10681 20033 10687
rect 20007 10649 20033 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 14239 10513 14265 10519
rect 14239 10481 14265 10487
rect 13959 10457 13985 10463
rect 8521 10431 8527 10457
rect 8553 10431 8559 10457
rect 13959 10425 13985 10431
rect 14631 10457 14657 10463
rect 14631 10425 14657 10431
rect 6231 10401 6257 10407
rect 13791 10401 13817 10407
rect 7233 10375 7239 10401
rect 7265 10375 7271 10401
rect 7513 10375 7519 10401
rect 7545 10375 7551 10401
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 10929 10375 10935 10401
rect 10961 10375 10967 10401
rect 6231 10369 6257 10375
rect 13791 10369 13817 10375
rect 13847 10401 13873 10407
rect 13847 10369 13873 10375
rect 14071 10401 14097 10407
rect 14071 10369 14097 10375
rect 7071 10345 7097 10351
rect 14183 10345 14209 10351
rect 11825 10319 11831 10345
rect 11857 10319 11863 10345
rect 7071 10313 7097 10319
rect 14183 10313 14209 10319
rect 14239 10345 14265 10351
rect 14239 10313 14265 10319
rect 6063 10289 6089 10295
rect 7401 10263 7407 10289
rect 7433 10263 7439 10289
rect 6063 10257 6089 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 11551 10121 11577 10127
rect 11551 10089 11577 10095
rect 12167 10121 12193 10127
rect 12167 10089 12193 10095
rect 8079 10065 8105 10071
rect 11775 10065 11801 10071
rect 5833 10039 5839 10065
rect 5865 10039 5871 10065
rect 7849 10039 7855 10065
rect 7881 10039 7887 10065
rect 8409 10039 8415 10065
rect 8441 10039 8447 10065
rect 8801 10039 8807 10065
rect 8833 10039 8839 10065
rect 10425 10039 10431 10065
rect 10457 10039 10463 10065
rect 11041 10039 11047 10065
rect 11073 10039 11079 10065
rect 8079 10033 8105 10039
rect 11775 10033 11801 10039
rect 12279 10065 12305 10071
rect 13455 10065 13481 10071
rect 12609 10039 12615 10065
rect 12641 10039 12647 10065
rect 12279 10033 12305 10039
rect 13455 10033 13481 10039
rect 13847 10065 13873 10071
rect 13847 10033 13873 10039
rect 7687 10009 7713 10015
rect 8639 10009 8665 10015
rect 12335 10009 12361 10015
rect 13623 10009 13649 10015
rect 5497 9983 5503 10009
rect 5529 9983 5535 10009
rect 7289 9983 7295 10009
rect 7321 9983 7327 10009
rect 8297 9983 8303 10009
rect 8329 9983 8335 10009
rect 8745 9983 8751 10009
rect 8777 9983 8783 10009
rect 8969 9983 8975 10009
rect 9001 9983 9007 10009
rect 9305 9983 9311 10009
rect 9337 9983 9343 10009
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 10929 9983 10935 10009
rect 10961 9983 10967 10009
rect 12721 9983 12727 10009
rect 12753 9983 12759 10009
rect 13225 9983 13231 10009
rect 13257 9983 13263 10009
rect 13337 9983 13343 10009
rect 13369 9983 13375 10009
rect 7687 9977 7713 9983
rect 8639 9977 8665 9983
rect 12335 9977 12361 9983
rect 13623 9977 13649 9983
rect 13735 10009 13761 10015
rect 13735 9977 13761 9983
rect 7519 9953 7545 9959
rect 6897 9927 6903 9953
rect 6929 9927 6935 9953
rect 7519 9921 7545 9927
rect 8023 9953 8049 9959
rect 13287 9953 13313 9959
rect 10761 9927 10767 9953
rect 10793 9927 10799 9953
rect 11993 9927 11999 9953
rect 12025 9927 12031 9953
rect 8023 9921 8049 9927
rect 13287 9921 13313 9927
rect 13679 9953 13705 9959
rect 13679 9921 13705 9927
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 10207 9729 10233 9735
rect 11153 9703 11159 9729
rect 11185 9703 11191 9729
rect 10207 9697 10233 9703
rect 20007 9673 20033 9679
rect 10313 9647 10319 9673
rect 10345 9647 10351 9673
rect 10985 9647 10991 9673
rect 11017 9647 11023 9673
rect 20007 9641 20033 9647
rect 7351 9617 7377 9623
rect 9255 9617 9281 9623
rect 8353 9591 8359 9617
rect 8385 9591 8391 9617
rect 8689 9591 8695 9617
rect 8721 9591 8727 9617
rect 9025 9591 9031 9617
rect 9057 9591 9063 9617
rect 7351 9585 7377 9591
rect 9255 9585 9281 9591
rect 9927 9617 9953 9623
rect 10369 9591 10375 9617
rect 10401 9591 10407 9617
rect 10929 9591 10935 9617
rect 10961 9591 10967 9617
rect 11097 9591 11103 9617
rect 11129 9591 11135 9617
rect 11825 9591 11831 9617
rect 11857 9591 11863 9617
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 9927 9585 9953 9591
rect 7519 9561 7545 9567
rect 9585 9535 9591 9561
rect 9617 9535 9623 9561
rect 9865 9535 9871 9561
rect 9897 9535 9903 9561
rect 13673 9535 13679 9561
rect 13705 9535 13711 9561
rect 7519 9529 7545 9535
rect 7015 9505 7041 9511
rect 7015 9473 7041 9479
rect 7407 9505 7433 9511
rect 8465 9479 8471 9505
rect 8497 9479 8503 9505
rect 8801 9479 8807 9505
rect 8833 9479 8839 9505
rect 9697 9479 9703 9505
rect 9729 9479 9735 9505
rect 7407 9473 7433 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 11103 9337 11129 9343
rect 11103 9305 11129 9311
rect 11663 9337 11689 9343
rect 11663 9305 11689 9311
rect 11775 9337 11801 9343
rect 12777 9311 12783 9337
rect 12809 9311 12815 9337
rect 11775 9305 11801 9311
rect 8751 9281 8777 9287
rect 12111 9281 12137 9287
rect 13511 9281 13537 9287
rect 9529 9255 9535 9281
rect 9561 9255 9567 9281
rect 10537 9255 10543 9281
rect 10569 9255 10575 9281
rect 13113 9255 13119 9281
rect 13145 9255 13151 9281
rect 8751 9249 8777 9255
rect 12111 9249 12137 9255
rect 13511 9249 13537 9255
rect 7295 9225 7321 9231
rect 5609 9199 5615 9225
rect 5641 9199 5647 9225
rect 6001 9199 6007 9225
rect 6033 9199 6039 9225
rect 7295 9193 7321 9199
rect 9255 9225 9281 9231
rect 11495 9225 11521 9231
rect 9473 9199 9479 9225
rect 9505 9199 9511 9225
rect 10033 9199 10039 9225
rect 10065 9199 10071 9225
rect 10257 9199 10263 9225
rect 10289 9199 10295 9225
rect 10761 9199 10767 9225
rect 10793 9199 10799 9225
rect 9255 9193 9281 9199
rect 11495 9193 11521 9199
rect 11943 9225 11969 9231
rect 11943 9193 11969 9199
rect 12615 9225 12641 9231
rect 13001 9199 13007 9225
rect 13033 9199 13039 9225
rect 13337 9199 13343 9225
rect 13369 9199 13375 9225
rect 13673 9199 13679 9225
rect 13705 9199 13711 9225
rect 12615 9193 12641 9199
rect 8807 9169 8833 9175
rect 7065 9143 7071 9169
rect 7097 9143 7103 9169
rect 8807 9137 8833 9143
rect 8975 9169 9001 9175
rect 10935 9169 10961 9175
rect 13455 9169 13481 9175
rect 9585 9143 9591 9169
rect 9617 9143 9623 9169
rect 10481 9143 10487 9169
rect 10513 9143 10519 9169
rect 10817 9143 10823 9169
rect 10849 9143 10855 9169
rect 11321 9143 11327 9169
rect 11353 9143 11359 9169
rect 11713 9143 11719 9169
rect 11745 9143 11751 9169
rect 14065 9143 14071 9169
rect 14097 9143 14103 9169
rect 15129 9143 15135 9169
rect 15161 9143 15167 9169
rect 8975 9137 9001 9143
rect 10935 9137 10961 9143
rect 13455 9137 13481 9143
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 9983 8945 10009 8951
rect 9983 8913 10009 8919
rect 10207 8945 10233 8951
rect 10207 8913 10233 8919
rect 10823 8945 10849 8951
rect 10823 8913 10849 8919
rect 12447 8945 12473 8951
rect 12447 8913 12473 8919
rect 14071 8945 14097 8951
rect 14071 8913 14097 8919
rect 9423 8889 9449 8895
rect 9423 8857 9449 8863
rect 10039 8889 10065 8895
rect 10039 8857 10065 8863
rect 10263 8889 10289 8895
rect 10263 8857 10289 8863
rect 10935 8889 10961 8895
rect 10935 8857 10961 8863
rect 11383 8889 11409 8895
rect 11383 8857 11409 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 8527 8833 8553 8839
rect 9143 8833 9169 8839
rect 11103 8833 11129 8839
rect 13959 8833 13985 8839
rect 14631 8833 14657 8839
rect 8745 8807 8751 8833
rect 8777 8807 8783 8833
rect 9473 8807 9479 8833
rect 9505 8807 9511 8833
rect 9697 8807 9703 8833
rect 9729 8807 9735 8833
rect 10369 8807 10375 8833
rect 10401 8807 10407 8833
rect 12441 8807 12447 8833
rect 12473 8807 12479 8833
rect 14177 8807 14183 8833
rect 14209 8807 14215 8833
rect 14737 8807 14743 8833
rect 14769 8807 14775 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 8527 8801 8553 8807
rect 9143 8801 9169 8807
rect 11103 8801 11129 8807
rect 13959 8801 13985 8807
rect 14631 8801 14657 8807
rect 9087 8777 9113 8783
rect 8857 8751 8863 8777
rect 8889 8751 8895 8777
rect 9087 8745 9113 8751
rect 12279 8777 12305 8783
rect 12279 8745 12305 8751
rect 14575 8777 14601 8783
rect 14575 8745 14601 8751
rect 8359 8721 8385 8727
rect 8359 8689 8385 8695
rect 8471 8721 8497 8727
rect 8471 8689 8497 8695
rect 8975 8721 9001 8727
rect 13511 8721 13537 8727
rect 10649 8695 10655 8721
rect 10681 8695 10687 8721
rect 8975 8689 9001 8695
rect 13511 8689 13537 8695
rect 14127 8721 14153 8727
rect 14127 8689 14153 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 8415 8553 8441 8559
rect 8415 8521 8441 8527
rect 8695 8553 8721 8559
rect 8695 8521 8721 8527
rect 10823 8553 10849 8559
rect 10823 8521 10849 8527
rect 13343 8553 13369 8559
rect 13343 8521 13369 8527
rect 9087 8497 9113 8503
rect 11215 8497 11241 8503
rect 7121 8471 7127 8497
rect 7153 8471 7159 8497
rect 9249 8471 9255 8497
rect 9281 8471 9287 8497
rect 10649 8471 10655 8497
rect 10681 8471 10687 8497
rect 9087 8465 9113 8471
rect 11215 8465 11241 8471
rect 12951 8497 12977 8503
rect 14177 8471 14183 8497
rect 14209 8471 14215 8497
rect 12951 8465 12977 8471
rect 9535 8441 9561 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 6785 8415 6791 8441
rect 6817 8415 6823 8441
rect 8801 8415 8807 8441
rect 8833 8415 8839 8441
rect 8969 8415 8975 8441
rect 9001 8415 9007 8441
rect 9535 8409 9561 8415
rect 11383 8441 11409 8447
rect 11383 8409 11409 8415
rect 11495 8441 11521 8447
rect 13623 8441 13649 8447
rect 13057 8415 13063 8441
rect 13089 8415 13095 8441
rect 13225 8415 13231 8441
rect 13257 8415 13263 8441
rect 13841 8415 13847 8441
rect 13873 8415 13879 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 11495 8409 11521 8415
rect 13623 8409 13649 8415
rect 11271 8385 11297 8391
rect 8185 8359 8191 8385
rect 8217 8359 8223 8385
rect 11271 8353 11297 8359
rect 12671 8385 12697 8391
rect 15241 8359 15247 8385
rect 15273 8359 15279 8385
rect 12671 8353 12697 8359
rect 967 8329 993 8335
rect 9423 8329 9449 8335
rect 20007 8329 20033 8335
rect 8801 8303 8807 8329
rect 8833 8303 8839 8329
rect 13225 8303 13231 8329
rect 13257 8303 13263 8329
rect 967 8297 993 8303
rect 9423 8297 9449 8303
rect 20007 8297 20033 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 10375 8161 10401 8167
rect 10375 8129 10401 8135
rect 13791 8161 13817 8167
rect 13791 8129 13817 8135
rect 13847 8105 13873 8111
rect 6729 8079 6735 8105
rect 6761 8079 6767 8105
rect 7793 8079 7799 8105
rect 7825 8079 7831 8105
rect 11265 8079 11271 8105
rect 11297 8079 11303 8105
rect 12329 8079 12335 8105
rect 12361 8079 12367 8105
rect 13847 8073 13873 8079
rect 8527 8049 8553 8055
rect 8185 8023 8191 8049
rect 8217 8023 8223 8049
rect 8353 8023 8359 8049
rect 8385 8023 8391 8049
rect 8527 8017 8553 8023
rect 8639 8049 8665 8055
rect 12503 8049 12529 8055
rect 10929 8023 10935 8049
rect 10961 8023 10967 8049
rect 8639 8017 8665 8023
rect 12503 8017 12529 8023
rect 12559 8049 12585 8055
rect 13001 8023 13007 8049
rect 13033 8023 13039 8049
rect 13953 8023 13959 8049
rect 13985 8023 13991 8049
rect 12559 8017 12585 8023
rect 10263 7993 10289 7999
rect 10263 7961 10289 7967
rect 8583 7937 8609 7943
rect 8583 7905 8609 7911
rect 10319 7937 10345 7943
rect 10319 7905 10345 7911
rect 12615 7937 12641 7943
rect 12615 7905 12641 7911
rect 12727 7937 12753 7943
rect 13113 7911 13119 7937
rect 13145 7911 13151 7937
rect 12727 7905 12753 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8303 7769 8329 7775
rect 8303 7737 8329 7743
rect 11887 7769 11913 7775
rect 11887 7737 11913 7743
rect 12839 7769 12865 7775
rect 12839 7737 12865 7743
rect 9255 7713 9281 7719
rect 12665 7687 12671 7713
rect 12697 7687 12703 7713
rect 13449 7687 13455 7713
rect 13481 7687 13487 7713
rect 9255 7681 9281 7687
rect 8807 7657 8833 7663
rect 8807 7625 8833 7631
rect 8919 7657 8945 7663
rect 8919 7625 8945 7631
rect 9087 7657 9113 7663
rect 9087 7625 9113 7631
rect 9143 7657 9169 7663
rect 9143 7625 9169 7631
rect 9311 7657 9337 7663
rect 9311 7625 9337 7631
rect 11999 7657 12025 7663
rect 11999 7625 12025 7631
rect 12223 7657 12249 7663
rect 14743 7657 14769 7663
rect 13057 7631 13063 7657
rect 13089 7631 13095 7657
rect 12223 7625 12249 7631
rect 14743 7625 14769 7631
rect 8975 7601 9001 7607
rect 8975 7569 9001 7575
rect 11943 7601 11969 7607
rect 14513 7575 14519 7601
rect 14545 7575 14551 7601
rect 11943 7569 11969 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9423 7377 9449 7383
rect 9423 7345 9449 7351
rect 8129 7295 8135 7321
rect 8161 7295 8167 7321
rect 9193 7295 9199 7321
rect 9225 7295 9231 7321
rect 9479 7265 9505 7271
rect 7793 7239 7799 7265
rect 7825 7239 7831 7265
rect 9479 7233 9505 7239
rect 9703 7265 9729 7271
rect 9703 7233 9729 7239
rect 10263 7265 10289 7271
rect 10263 7233 10289 7239
rect 10375 7265 10401 7271
rect 10375 7233 10401 7239
rect 10655 7265 10681 7271
rect 10655 7233 10681 7239
rect 10991 7265 11017 7271
rect 10991 7233 11017 7239
rect 12559 7265 12585 7271
rect 12559 7233 12585 7239
rect 12671 7265 12697 7271
rect 12671 7233 12697 7239
rect 13119 7265 13145 7271
rect 13119 7233 13145 7239
rect 10095 7209 10121 7215
rect 10095 7177 10121 7183
rect 10767 7209 10793 7215
rect 10767 7177 10793 7183
rect 12839 7209 12865 7215
rect 12839 7177 12865 7183
rect 12951 7209 12977 7215
rect 12951 7177 12977 7183
rect 9423 7153 9449 7159
rect 9423 7121 9449 7127
rect 10207 7153 10233 7159
rect 10207 7121 10233 7127
rect 10823 7153 10849 7159
rect 10823 7121 10849 7127
rect 12783 7153 12809 7159
rect 12783 7121 12809 7127
rect 13063 7153 13089 7159
rect 13063 7121 13089 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 11999 6985 12025 6991
rect 11999 6953 12025 6959
rect 14295 6985 14321 6991
rect 14295 6953 14321 6959
rect 8807 6929 8833 6935
rect 8807 6897 8833 6903
rect 8975 6929 9001 6935
rect 8975 6897 9001 6903
rect 9983 6929 10009 6935
rect 9983 6897 10009 6903
rect 10095 6929 10121 6935
rect 10095 6897 10121 6903
rect 10151 6929 10177 6935
rect 10705 6903 10711 6929
rect 10737 6903 10743 6929
rect 13001 6903 13007 6929
rect 13033 6903 13039 6929
rect 10151 6897 10177 6903
rect 9031 6873 9057 6879
rect 10313 6847 10319 6873
rect 10345 6847 10351 6873
rect 12609 6847 12615 6873
rect 12641 6847 12647 6873
rect 9031 6841 9057 6847
rect 8863 6817 8889 6823
rect 11769 6791 11775 6817
rect 11801 6791 11807 6817
rect 14065 6791 14071 6817
rect 14097 6791 14103 6817
rect 8863 6785 8889 6791
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 9423 6537 9449 6543
rect 8129 6511 8135 6537
rect 8161 6511 8167 6537
rect 9193 6511 9199 6537
rect 9225 6511 9231 6537
rect 9423 6505 9449 6511
rect 7793 6455 7799 6481
rect 7825 6455 7831 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 9423 6201 9449 6207
rect 9423 6169 9449 6175
rect 9977 6119 9983 6145
rect 10009 6119 10015 6145
rect 9585 6063 9591 6089
rect 9617 6063 9623 6089
rect 11041 6007 11047 6033
rect 11073 6007 11079 6033
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 13007 2617 13033 2623
rect 13007 2585 13033 2591
rect 13953 2535 13959 2561
rect 13985 2535 13991 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9641 2143 9647 2169
rect 9673 2143 9679 2169
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 10039 2057 10065 2063
rect 10039 2025 10065 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 11215 1833 11241 1839
rect 11215 1801 11241 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 9025 1751 9031 1777
rect 9057 1751 9063 1777
rect 10873 1751 10879 1777
rect 10905 1751 10911 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 8807 18999 8833 19025
rect 10711 18999 10737 19025
rect 12279 18999 12305 19025
rect 3151 18943 3177 18969
rect 10487 18943 10513 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9199 18719 9225 18745
rect 10711 18719 10737 18745
rect 8695 18607 8721 18633
rect 10207 18607 10233 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9927 14239 9953 14265
rect 9983 14239 10009 14265
rect 10263 14239 10289 14265
rect 10319 14239 10345 14265
rect 9815 14183 9841 14209
rect 10431 14183 10457 14209
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8751 14015 8777 14041
rect 8807 13959 8833 13985
rect 7015 13903 7041 13929
rect 8639 13903 8665 13929
rect 9591 13903 9617 13929
rect 7351 13847 7377 13873
rect 8415 13847 8441 13873
rect 9087 13847 9113 13873
rect 9479 13847 9505 13873
rect 9983 13847 10009 13873
rect 11047 13847 11073 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 8191 13567 8217 13593
rect 8527 13567 8553 13593
rect 10375 13567 10401 13593
rect 10823 13567 10849 13593
rect 20007 13567 20033 13593
rect 6791 13511 6817 13537
rect 8639 13511 8665 13537
rect 8919 13511 8945 13537
rect 18831 13511 18857 13537
rect 7127 13455 7153 13481
rect 8471 13455 8497 13481
rect 8751 13455 8777 13481
rect 9311 13455 9337 13481
rect 10655 13455 10681 13481
rect 10767 13399 10793 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7631 13231 7657 13257
rect 8751 13231 8777 13257
rect 9591 13231 9617 13257
rect 10039 13231 10065 13257
rect 8023 13175 8049 13201
rect 8191 13175 8217 13201
rect 8975 13175 9001 13201
rect 9703 13175 9729 13201
rect 9815 13175 9841 13201
rect 10151 13175 10177 13201
rect 10263 13175 10289 13201
rect 10879 13175 10905 13201
rect 13063 13175 13089 13201
rect 7519 13119 7545 13145
rect 8303 13119 8329 13145
rect 9087 13119 9113 13145
rect 9535 13119 9561 13145
rect 9927 13119 9953 13145
rect 10543 13119 10569 13145
rect 12839 13119 12865 13145
rect 12951 13119 12977 13145
rect 18943 13119 18969 13145
rect 8079 13063 8105 13089
rect 11943 13063 11969 13089
rect 12223 13063 12249 13089
rect 13679 13063 13705 13089
rect 19951 13063 19977 13089
rect 7687 13007 7713 13033
rect 12895 13007 12921 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 967 12783 993 12809
rect 8303 12783 8329 12809
rect 10767 12783 10793 12809
rect 13511 12783 13537 12809
rect 20007 12783 20033 12809
rect 2143 12727 2169 12753
rect 10991 12727 11017 12753
rect 12111 12727 12137 12753
rect 14183 12727 14209 12753
rect 18831 12727 18857 12753
rect 8527 12671 8553 12697
rect 12447 12671 12473 12697
rect 13791 12671 13817 12697
rect 14295 12671 14321 12697
rect 8695 12615 8721 12641
rect 10711 12615 10737 12641
rect 10767 12615 10793 12641
rect 10879 12615 10905 12641
rect 13623 12615 13649 12641
rect 13735 12615 13761 12641
rect 14575 12615 14601 12641
rect 14743 12615 14769 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8191 12447 8217 12473
rect 9871 12447 9897 12473
rect 12783 12447 12809 12473
rect 8919 12391 8945 12417
rect 9927 12391 9953 12417
rect 13399 12391 13425 12417
rect 7967 12335 7993 12361
rect 8695 12335 8721 12361
rect 8807 12335 8833 12361
rect 10039 12335 10065 12361
rect 10151 12335 10177 12361
rect 13007 12335 13033 12361
rect 18831 12335 18857 12361
rect 6511 12279 6537 12305
rect 7575 12279 7601 12305
rect 8751 12279 8777 12305
rect 14519 12279 14545 12305
rect 14799 12279 14825 12305
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 7575 12055 7601 12081
rect 8191 11999 8217 12025
rect 9535 11999 9561 12025
rect 12671 11999 12697 12025
rect 13343 11999 13369 12025
rect 20007 11999 20033 12025
rect 7743 11943 7769 11969
rect 8135 11943 8161 11969
rect 8247 11943 8273 11969
rect 8359 11943 8385 11969
rect 8471 11943 8497 11969
rect 10095 11943 10121 11969
rect 11271 11943 11297 11969
rect 12783 11943 12809 11969
rect 12951 11943 12977 11969
rect 13175 11943 13201 11969
rect 13287 11943 13313 11969
rect 18831 11943 18857 11969
rect 7631 11887 7657 11913
rect 9479 11887 9505 11913
rect 9535 11887 9561 11913
rect 9591 11887 9617 11913
rect 11607 11887 11633 11913
rect 13399 11887 13425 11913
rect 9703 11831 9729 11857
rect 10151 11831 10177 11857
rect 10263 11831 10289 11857
rect 12895 11831 12921 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 8023 11663 8049 11689
rect 9367 11663 9393 11689
rect 10543 11663 10569 11689
rect 11775 11663 11801 11689
rect 12671 11663 12697 11689
rect 12951 11663 12977 11689
rect 7575 11607 7601 11633
rect 9143 11607 9169 11633
rect 9199 11607 9225 11633
rect 10095 11607 10121 11633
rect 10375 11607 10401 11633
rect 10655 11607 10681 11633
rect 12727 11607 12753 11633
rect 2143 11551 2169 11577
rect 7351 11551 7377 11577
rect 7743 11551 7769 11577
rect 7911 11551 7937 11577
rect 8247 11551 8273 11577
rect 9031 11551 9057 11577
rect 9535 11551 9561 11577
rect 9703 11551 9729 11577
rect 9927 11551 9953 11577
rect 10823 11551 10849 11577
rect 11551 11551 11577 11577
rect 11719 11551 11745 11577
rect 11887 11551 11913 11577
rect 12559 11551 12585 11577
rect 5895 11495 5921 11521
rect 6959 11495 6985 11521
rect 8135 11495 8161 11521
rect 967 11439 993 11465
rect 8023 11439 8049 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7407 11271 7433 11297
rect 7575 11271 7601 11297
rect 7967 11271 7993 11297
rect 13063 11271 13089 11297
rect 11383 11215 11409 11241
rect 20007 11215 20033 11241
rect 9479 11159 9505 11185
rect 9591 11159 9617 11185
rect 10655 11159 10681 11185
rect 12839 11159 12865 11185
rect 13119 11159 13145 11185
rect 13231 11159 13257 11185
rect 13287 11159 13313 11185
rect 18831 11159 18857 11185
rect 7911 11103 7937 11129
rect 9871 11103 9897 11129
rect 10767 11103 10793 11129
rect 11103 11103 11129 11129
rect 12447 11103 12473 11129
rect 13007 11103 13033 11129
rect 7463 11047 7489 11073
rect 7967 11047 7993 11073
rect 9367 11047 9393 11073
rect 10935 11047 10961 11073
rect 14295 11047 14321 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 9815 10879 9841 10905
rect 8415 10823 8441 10849
rect 9143 10823 9169 10849
rect 9759 10823 9785 10849
rect 11607 10823 11633 10849
rect 11999 10823 12025 10849
rect 13231 10823 13257 10849
rect 7183 10767 7209 10793
rect 7799 10767 7825 10793
rect 8191 10767 8217 10793
rect 8303 10767 8329 10793
rect 8919 10767 8945 10793
rect 9815 10767 9841 10793
rect 10487 10767 10513 10793
rect 11159 10767 11185 10793
rect 11775 10767 11801 10793
rect 12055 10767 12081 10793
rect 12839 10767 12865 10793
rect 14519 10767 14545 10793
rect 18831 10767 18857 10793
rect 6847 10711 6873 10737
rect 7295 10711 7321 10737
rect 7575 10711 7601 10737
rect 8359 10711 8385 10737
rect 14295 10711 14321 10737
rect 14855 10711 14881 10737
rect 15919 10711 15945 10737
rect 11999 10655 12025 10681
rect 20007 10655 20033 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 14239 10487 14265 10513
rect 8527 10431 8553 10457
rect 13959 10431 13985 10457
rect 14631 10431 14657 10457
rect 6231 10375 6257 10401
rect 7239 10375 7265 10401
rect 7519 10375 7545 10401
rect 10039 10375 10065 10401
rect 10935 10375 10961 10401
rect 13791 10375 13817 10401
rect 13847 10375 13873 10401
rect 14071 10375 14097 10401
rect 7071 10319 7097 10345
rect 11831 10319 11857 10345
rect 14183 10319 14209 10345
rect 14239 10319 14265 10345
rect 6063 10263 6089 10289
rect 7407 10263 7433 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 11551 10095 11577 10121
rect 12167 10095 12193 10121
rect 5839 10039 5865 10065
rect 7855 10039 7881 10065
rect 8079 10039 8105 10065
rect 8415 10039 8441 10065
rect 8807 10039 8833 10065
rect 10431 10039 10457 10065
rect 11047 10039 11073 10065
rect 11775 10039 11801 10065
rect 12279 10039 12305 10065
rect 12615 10039 12641 10065
rect 13455 10039 13481 10065
rect 13847 10039 13873 10065
rect 5503 9983 5529 10009
rect 7295 9983 7321 10009
rect 7687 9983 7713 10009
rect 8303 9983 8329 10009
rect 8639 9983 8665 10009
rect 8751 9983 8777 10009
rect 8975 9983 9001 10009
rect 9311 9983 9337 10009
rect 9703 9983 9729 10009
rect 10935 9983 10961 10009
rect 12335 9983 12361 10009
rect 12727 9983 12753 10009
rect 13231 9983 13257 10009
rect 13343 9983 13369 10009
rect 13623 9983 13649 10009
rect 13735 9983 13761 10009
rect 6903 9927 6929 9953
rect 7519 9927 7545 9953
rect 8023 9927 8049 9953
rect 10767 9927 10793 9953
rect 11999 9927 12025 9953
rect 13287 9927 13313 9953
rect 13679 9927 13705 9953
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 10207 9703 10233 9729
rect 11159 9703 11185 9729
rect 10319 9647 10345 9673
rect 10991 9647 11017 9673
rect 20007 9647 20033 9673
rect 7351 9591 7377 9617
rect 8359 9591 8385 9617
rect 8695 9591 8721 9617
rect 9031 9591 9057 9617
rect 9255 9591 9281 9617
rect 9927 9591 9953 9617
rect 10375 9591 10401 9617
rect 10935 9591 10961 9617
rect 11103 9591 11129 9617
rect 11831 9591 11857 9617
rect 18831 9591 18857 9617
rect 7519 9535 7545 9561
rect 9591 9535 9617 9561
rect 9871 9535 9897 9561
rect 13679 9535 13705 9561
rect 7015 9479 7041 9505
rect 7407 9479 7433 9505
rect 8471 9479 8497 9505
rect 8807 9479 8833 9505
rect 9703 9479 9729 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 11103 9311 11129 9337
rect 11663 9311 11689 9337
rect 11775 9311 11801 9337
rect 12783 9311 12809 9337
rect 8751 9255 8777 9281
rect 9535 9255 9561 9281
rect 10543 9255 10569 9281
rect 12111 9255 12137 9281
rect 13119 9255 13145 9281
rect 13511 9255 13537 9281
rect 5615 9199 5641 9225
rect 6007 9199 6033 9225
rect 7295 9199 7321 9225
rect 9255 9199 9281 9225
rect 9479 9199 9505 9225
rect 10039 9199 10065 9225
rect 10263 9199 10289 9225
rect 10767 9199 10793 9225
rect 11495 9199 11521 9225
rect 11943 9199 11969 9225
rect 12615 9199 12641 9225
rect 13007 9199 13033 9225
rect 13343 9199 13369 9225
rect 13679 9199 13705 9225
rect 7071 9143 7097 9169
rect 8807 9143 8833 9169
rect 8975 9143 9001 9169
rect 9591 9143 9617 9169
rect 10487 9143 10513 9169
rect 10823 9143 10849 9169
rect 10935 9143 10961 9169
rect 11327 9143 11353 9169
rect 11719 9143 11745 9169
rect 13455 9143 13481 9169
rect 14071 9143 14097 9169
rect 15135 9143 15161 9169
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 9983 8919 10009 8945
rect 10207 8919 10233 8945
rect 10823 8919 10849 8945
rect 12447 8919 12473 8945
rect 14071 8919 14097 8945
rect 9423 8863 9449 8889
rect 10039 8863 10065 8889
rect 10263 8863 10289 8889
rect 10935 8863 10961 8889
rect 11383 8863 11409 8889
rect 20007 8863 20033 8889
rect 8527 8807 8553 8833
rect 8751 8807 8777 8833
rect 9143 8807 9169 8833
rect 9479 8807 9505 8833
rect 9703 8807 9729 8833
rect 10375 8807 10401 8833
rect 11103 8807 11129 8833
rect 12447 8807 12473 8833
rect 13959 8807 13985 8833
rect 14183 8807 14209 8833
rect 14631 8807 14657 8833
rect 14743 8807 14769 8833
rect 18831 8807 18857 8833
rect 8863 8751 8889 8777
rect 9087 8751 9113 8777
rect 12279 8751 12305 8777
rect 14575 8751 14601 8777
rect 8359 8695 8385 8721
rect 8471 8695 8497 8721
rect 8975 8695 9001 8721
rect 10655 8695 10681 8721
rect 13511 8695 13537 8721
rect 14127 8695 14153 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 8415 8527 8441 8553
rect 8695 8527 8721 8553
rect 10823 8527 10849 8553
rect 13343 8527 13369 8553
rect 7127 8471 7153 8497
rect 9087 8471 9113 8497
rect 9255 8471 9281 8497
rect 10655 8471 10681 8497
rect 11215 8471 11241 8497
rect 12951 8471 12977 8497
rect 14183 8471 14209 8497
rect 2143 8415 2169 8441
rect 6791 8415 6817 8441
rect 8807 8415 8833 8441
rect 8975 8415 9001 8441
rect 9535 8415 9561 8441
rect 11383 8415 11409 8441
rect 11495 8415 11521 8441
rect 13063 8415 13089 8441
rect 13231 8415 13257 8441
rect 13623 8415 13649 8441
rect 13847 8415 13873 8441
rect 18831 8415 18857 8441
rect 8191 8359 8217 8385
rect 11271 8359 11297 8385
rect 12671 8359 12697 8385
rect 15247 8359 15273 8385
rect 967 8303 993 8329
rect 8807 8303 8833 8329
rect 9423 8303 9449 8329
rect 13231 8303 13257 8329
rect 20007 8303 20033 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 10375 8135 10401 8161
rect 13791 8135 13817 8161
rect 6735 8079 6761 8105
rect 7799 8079 7825 8105
rect 11271 8079 11297 8105
rect 12335 8079 12361 8105
rect 13847 8079 13873 8105
rect 8191 8023 8217 8049
rect 8359 8023 8385 8049
rect 8527 8023 8553 8049
rect 8639 8023 8665 8049
rect 10935 8023 10961 8049
rect 12503 8023 12529 8049
rect 12559 8023 12585 8049
rect 13007 8023 13033 8049
rect 13959 8023 13985 8049
rect 10263 7967 10289 7993
rect 8583 7911 8609 7937
rect 10319 7911 10345 7937
rect 12615 7911 12641 7937
rect 12727 7911 12753 7937
rect 13119 7911 13145 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8303 7743 8329 7769
rect 11887 7743 11913 7769
rect 12839 7743 12865 7769
rect 9255 7687 9281 7713
rect 12671 7687 12697 7713
rect 13455 7687 13481 7713
rect 8807 7631 8833 7657
rect 8919 7631 8945 7657
rect 9087 7631 9113 7657
rect 9143 7631 9169 7657
rect 9311 7631 9337 7657
rect 11999 7631 12025 7657
rect 12223 7631 12249 7657
rect 13063 7631 13089 7657
rect 14743 7631 14769 7657
rect 8975 7575 9001 7601
rect 11943 7575 11969 7601
rect 14519 7575 14545 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9423 7351 9449 7377
rect 8135 7295 8161 7321
rect 9199 7295 9225 7321
rect 7799 7239 7825 7265
rect 9479 7239 9505 7265
rect 9703 7239 9729 7265
rect 10263 7239 10289 7265
rect 10375 7239 10401 7265
rect 10655 7239 10681 7265
rect 10991 7239 11017 7265
rect 12559 7239 12585 7265
rect 12671 7239 12697 7265
rect 13119 7239 13145 7265
rect 10095 7183 10121 7209
rect 10767 7183 10793 7209
rect 12839 7183 12865 7209
rect 12951 7183 12977 7209
rect 9423 7127 9449 7153
rect 10207 7127 10233 7153
rect 10823 7127 10849 7153
rect 12783 7127 12809 7153
rect 13063 7127 13089 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 11999 6959 12025 6985
rect 14295 6959 14321 6985
rect 8807 6903 8833 6929
rect 8975 6903 9001 6929
rect 9983 6903 10009 6929
rect 10095 6903 10121 6929
rect 10151 6903 10177 6929
rect 10711 6903 10737 6929
rect 13007 6903 13033 6929
rect 9031 6847 9057 6873
rect 10319 6847 10345 6873
rect 12615 6847 12641 6873
rect 8863 6791 8889 6817
rect 11775 6791 11801 6817
rect 14071 6791 14097 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8135 6511 8161 6537
rect 9199 6511 9225 6537
rect 9423 6511 9449 6537
rect 7799 6455 7825 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 9423 6175 9449 6201
rect 9983 6119 10009 6145
rect 9591 6063 9617 6089
rect 11047 6007 11073 6033
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 13007 2591 13033 2617
rect 13959 2535 13985 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9647 2143 9673 2169
rect 12615 2143 12641 2169
rect 10039 2031 10065 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 11215 1807 11241 1833
rect 12783 1807 12809 1833
rect 9031 1751 9057 1777
rect 10879 1751 10905 1777
rect 12279 1751 12305 1777
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 3024 20600 3080 21000
rect 8064 20600 8120 21000
rect 8736 20600 8792 21000
rect 10080 20600 10136 21000
rect 10416 20600 10472 21000
rect 10752 20600 10808 21000
rect 11760 20600 11816 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 3038 18970 3066 20600
rect 3150 18970 3178 18975
rect 3038 18969 3178 18970
rect 3038 18943 3151 18969
rect 3177 18943 3178 18969
rect 3038 18942 3178 18943
rect 3150 18937 3178 18942
rect 8078 18746 8106 20600
rect 8750 19138 8778 20600
rect 8750 19105 8778 19110
rect 9310 19138 9338 19143
rect 9310 19091 9338 19110
rect 8078 18713 8106 18718
rect 8806 19025 8834 19031
rect 8806 18999 8807 19025
rect 8833 18999 8834 19025
rect 8694 18633 8722 18639
rect 8694 18607 8695 18633
rect 8721 18607 8722 18633
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 8190 14210 8218 14215
rect 7014 13929 7042 13935
rect 7014 13903 7015 13929
rect 7041 13903 7042 13929
rect 2086 13818 2114 13823
rect 966 12809 994 12815
rect 966 12783 967 12809
rect 993 12783 994 12809
rect 966 12474 994 12783
rect 966 12441 994 12446
rect 966 11466 994 11471
rect 966 11419 994 11438
rect 2086 10402 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 6790 13538 6818 13543
rect 7014 13538 7042 13903
rect 7350 13874 7378 13879
rect 7350 13827 7378 13846
rect 6790 13537 7042 13538
rect 6790 13511 6791 13537
rect 6817 13511 7042 13537
rect 6790 13510 7042 13511
rect 6790 13505 6818 13510
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2142 12754 2170 12759
rect 2142 12707 2170 12726
rect 6510 12754 6538 12759
rect 6510 12305 6538 12726
rect 7014 12642 7042 13510
rect 8190 13593 8218 14182
rect 8694 14210 8722 18607
rect 8806 15974 8834 18999
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9198 18746 9226 18751
rect 9198 18699 9226 18718
rect 10094 18746 10122 20600
rect 10430 18970 10458 20600
rect 10766 19138 10794 20600
rect 10766 19105 10794 19110
rect 11214 19138 11242 19143
rect 11214 19091 11242 19110
rect 11774 19138 11802 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 11774 19105 11802 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 10710 19026 10738 19031
rect 10654 19025 10738 19026
rect 10654 18999 10711 19025
rect 10737 18999 10738 19025
rect 10654 18998 10738 18999
rect 10486 18970 10514 18975
rect 10430 18969 10514 18970
rect 10430 18943 10487 18969
rect 10513 18943 10514 18969
rect 10430 18942 10514 18943
rect 10486 18937 10514 18942
rect 10094 18713 10122 18718
rect 10206 18633 10234 18639
rect 10206 18607 10207 18633
rect 10233 18607 10234 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 10206 15974 10234 18607
rect 10654 15974 10682 18998
rect 10710 18993 10738 18998
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 10710 18746 10738 18751
rect 10710 18699 10738 18718
rect 12278 15974 12306 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 8694 14177 8722 14182
rect 8750 15946 8834 15974
rect 10094 15946 10234 15974
rect 10318 15946 10682 15974
rect 11942 15946 12306 15974
rect 8750 14042 8778 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 10094 14378 10122 15946
rect 9926 14350 10122 14378
rect 9926 14266 9954 14350
rect 9926 14219 9954 14238
rect 9982 14266 10010 14271
rect 10262 14266 10290 14271
rect 9982 14265 10290 14266
rect 9982 14239 9983 14265
rect 10009 14239 10263 14265
rect 10289 14239 10290 14265
rect 9982 14238 10290 14239
rect 8414 14041 8778 14042
rect 8414 14015 8751 14041
rect 8777 14015 8778 14041
rect 8414 14014 8778 14015
rect 8414 13873 8442 14014
rect 8750 14009 8778 14014
rect 8806 14210 8834 14215
rect 9814 14210 9842 14215
rect 8806 13985 8834 14182
rect 8806 13959 8807 13985
rect 8833 13959 8834 13985
rect 8638 13929 8666 13935
rect 8638 13903 8639 13929
rect 8665 13903 8666 13929
rect 8414 13847 8415 13873
rect 8441 13847 8442 13873
rect 8414 13841 8442 13847
rect 8526 13874 8554 13879
rect 8190 13567 8191 13593
rect 8217 13567 8218 13593
rect 7126 13481 7154 13487
rect 7126 13455 7127 13481
rect 7153 13455 7154 13481
rect 7126 13370 7154 13455
rect 8022 13426 8050 13431
rect 7126 13337 7154 13342
rect 7574 13370 7602 13375
rect 7602 13342 7658 13370
rect 7574 13337 7602 13342
rect 7630 13257 7658 13342
rect 7630 13231 7631 13257
rect 7657 13231 7658 13257
rect 7630 13225 7658 13231
rect 8022 13201 8050 13398
rect 8022 13175 8023 13201
rect 8049 13175 8050 13201
rect 8022 13169 8050 13175
rect 8190 13201 8218 13567
rect 8526 13593 8554 13846
rect 8526 13567 8527 13593
rect 8553 13567 8554 13593
rect 8526 13561 8554 13567
rect 8638 13537 8666 13903
rect 8638 13511 8639 13537
rect 8665 13511 8666 13537
rect 8638 13505 8666 13511
rect 8190 13175 8191 13201
rect 8217 13175 8218 13201
rect 8190 13169 8218 13175
rect 8470 13481 8498 13487
rect 8470 13455 8471 13481
rect 8497 13455 8498 13481
rect 7518 13146 7546 13151
rect 7630 13146 7658 13151
rect 7518 13145 7630 13146
rect 7518 13119 7519 13145
rect 7545 13119 7630 13145
rect 7518 13118 7630 13119
rect 7518 13113 7546 13118
rect 7014 12609 7042 12614
rect 6510 12279 6511 12305
rect 6537 12279 6538 12305
rect 6510 12250 6538 12279
rect 6510 12217 6538 12222
rect 7574 12305 7602 12311
rect 7574 12279 7575 12305
rect 7601 12279 7602 12305
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 7574 12081 7602 12279
rect 7574 12055 7575 12081
rect 7601 12055 7602 12081
rect 7574 12049 7602 12055
rect 7630 11913 7658 13118
rect 8302 13146 8330 13151
rect 8302 13145 8386 13146
rect 8302 13119 8303 13145
rect 8329 13119 8386 13145
rect 8302 13118 8386 13119
rect 8302 13113 8330 13118
rect 8078 13089 8106 13095
rect 8078 13063 8079 13089
rect 8105 13063 8106 13089
rect 7686 13034 7714 13039
rect 8078 13034 8106 13063
rect 7686 13033 8106 13034
rect 7686 13007 7687 13033
rect 7713 13007 8106 13033
rect 7686 13006 8106 13007
rect 7686 13001 7714 13006
rect 8302 12810 8330 12815
rect 8190 12782 8302 12810
rect 7966 12642 7994 12647
rect 7966 12474 7994 12614
rect 8190 12474 8218 12782
rect 8302 12763 8330 12782
rect 8358 12698 8386 13118
rect 8302 12670 8386 12698
rect 7966 12473 8218 12474
rect 7966 12447 8191 12473
rect 8217 12447 8218 12473
rect 7966 12446 8218 12447
rect 7966 12361 7994 12446
rect 8190 12441 8218 12446
rect 8246 12642 8274 12647
rect 8246 12362 8274 12614
rect 7966 12335 7967 12361
rect 7993 12335 7994 12361
rect 7742 11970 7770 11975
rect 7742 11923 7770 11942
rect 7630 11887 7631 11913
rect 7657 11887 7658 11913
rect 7630 11746 7658 11887
rect 7966 11802 7994 12335
rect 8134 12334 8274 12362
rect 8134 11970 8162 12334
rect 8246 12250 8274 12255
rect 7966 11769 7994 11774
rect 8078 11969 8162 11970
rect 8078 11943 8135 11969
rect 8161 11943 8162 11969
rect 8078 11942 8162 11943
rect 7518 11718 7658 11746
rect 2142 11578 2170 11583
rect 2142 11531 2170 11550
rect 5894 11578 5922 11583
rect 5894 11521 5922 11550
rect 7350 11577 7378 11583
rect 7350 11551 7351 11577
rect 7377 11551 7378 11577
rect 5894 11495 5895 11521
rect 5921 11495 5922 11521
rect 5894 11489 5922 11495
rect 6958 11522 6986 11527
rect 7350 11522 7378 11551
rect 6958 11521 7266 11522
rect 6958 11495 6959 11521
rect 6985 11495 7266 11521
rect 6958 11494 7266 11495
rect 6958 11489 6986 11494
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 7238 11354 7266 11494
rect 7350 11489 7378 11494
rect 7238 11326 7434 11354
rect 7406 11297 7434 11326
rect 7406 11271 7407 11297
rect 7433 11271 7434 11297
rect 7406 11265 7434 11271
rect 7462 11074 7490 11079
rect 7518 11074 7546 11718
rect 8022 11690 8050 11695
rect 7630 11689 8050 11690
rect 7630 11663 8023 11689
rect 8049 11663 8050 11689
rect 7630 11662 8050 11663
rect 7574 11634 7602 11639
rect 7574 11522 7602 11606
rect 7574 11489 7602 11494
rect 7574 11298 7602 11303
rect 7630 11298 7658 11662
rect 8022 11657 8050 11662
rect 7742 11578 7770 11583
rect 7742 11531 7770 11550
rect 7910 11578 7938 11583
rect 7910 11531 7938 11550
rect 8078 11578 8106 11942
rect 8134 11937 8162 11942
rect 8190 12025 8218 12031
rect 8190 11999 8191 12025
rect 8217 11999 8218 12025
rect 8190 11970 8218 11999
rect 8190 11937 8218 11942
rect 8246 11969 8274 12222
rect 8246 11943 8247 11969
rect 8273 11943 8274 11969
rect 8246 11937 8274 11943
rect 8302 11746 8330 12670
rect 8470 12530 8498 13455
rect 8750 13481 8778 13487
rect 8750 13455 8751 13481
rect 8777 13455 8778 13481
rect 8750 13454 8778 13455
rect 8526 13426 8554 13431
rect 8526 12697 8554 13398
rect 8694 13426 8778 13454
rect 8806 13426 8834 13959
rect 9702 14209 9842 14210
rect 9702 14183 9815 14209
rect 9841 14183 9842 14209
rect 9702 14182 9842 14183
rect 9590 13929 9618 13935
rect 9590 13903 9591 13929
rect 9617 13903 9618 13929
rect 9086 13874 9114 13879
rect 8918 13538 8946 13543
rect 9086 13538 9114 13846
rect 9478 13874 9506 13879
rect 9590 13874 9618 13903
rect 9506 13846 9618 13874
rect 9478 13827 9506 13846
rect 8918 13537 9114 13538
rect 8918 13511 8919 13537
rect 8945 13511 9114 13537
rect 8918 13510 9114 13511
rect 8918 13454 8946 13510
rect 8694 13202 8722 13426
rect 8806 13393 8834 13398
rect 8862 13426 8946 13454
rect 9310 13482 9338 13487
rect 9310 13481 9618 13482
rect 9310 13455 9311 13481
rect 9337 13455 9618 13481
rect 9310 13454 9618 13455
rect 9310 13449 9338 13454
rect 8862 13314 8890 13426
rect 8694 13169 8722 13174
rect 8750 13286 8890 13314
rect 8750 13257 8778 13286
rect 8750 13231 8751 13257
rect 8777 13231 8778 13257
rect 8750 12810 8778 13231
rect 9590 13257 9618 13454
rect 9590 13231 9591 13257
rect 9617 13231 9618 13257
rect 9590 13225 9618 13231
rect 8974 13202 9002 13207
rect 8974 13155 9002 13174
rect 9702 13201 9730 14182
rect 9814 14177 9842 14182
rect 9982 14210 10010 14238
rect 10262 14233 10290 14238
rect 10318 14266 10346 15946
rect 10318 14219 10346 14238
rect 11046 14266 11074 14271
rect 9982 14177 10010 14182
rect 10374 14210 10402 14215
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9982 13873 10010 13879
rect 9982 13847 9983 13873
rect 10009 13847 10010 13873
rect 9982 13426 10010 13847
rect 10374 13593 10402 14182
rect 10374 13567 10375 13593
rect 10401 13567 10402 13593
rect 10374 13561 10402 13567
rect 10430 14209 10458 14215
rect 10430 14183 10431 14209
rect 10457 14183 10458 14209
rect 10430 13482 10458 14183
rect 11046 13873 11074 14238
rect 11046 13847 11047 13873
rect 11073 13847 11074 13873
rect 11046 13841 11074 13847
rect 10822 13594 10850 13599
rect 10822 13593 10906 13594
rect 10822 13567 10823 13593
rect 10849 13567 10906 13593
rect 10822 13566 10906 13567
rect 10822 13561 10850 13566
rect 10150 13454 10458 13482
rect 10654 13481 10682 13487
rect 10654 13455 10655 13481
rect 10681 13455 10682 13481
rect 9982 13398 10122 13426
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10038 13258 10066 13263
rect 10094 13258 10122 13398
rect 10038 13257 10122 13258
rect 10038 13231 10039 13257
rect 10065 13231 10122 13257
rect 10038 13230 10122 13231
rect 10038 13225 10066 13230
rect 9702 13175 9703 13201
rect 9729 13175 9730 13201
rect 9702 13169 9730 13175
rect 9814 13202 9842 13207
rect 9814 13155 9842 13174
rect 10150 13201 10178 13454
rect 10150 13175 10151 13201
rect 10177 13175 10178 13201
rect 10150 13169 10178 13175
rect 10262 13202 10290 13207
rect 10262 13155 10290 13174
rect 10654 13202 10682 13455
rect 10654 13169 10682 13174
rect 10766 13425 10794 13431
rect 10766 13399 10767 13425
rect 10793 13399 10794 13425
rect 9086 13146 9114 13151
rect 9086 13099 9114 13118
rect 9534 13145 9562 13151
rect 9534 13119 9535 13145
rect 9561 13119 9562 13145
rect 8750 12777 8778 12782
rect 8526 12671 8527 12697
rect 8553 12671 8554 12697
rect 8526 12665 8554 12671
rect 8694 12642 8722 12647
rect 8694 12595 8722 12614
rect 9366 12642 9394 12647
rect 8470 12502 8778 12530
rect 8358 12362 8386 12367
rect 8358 11969 8386 12334
rect 8694 12362 8722 12367
rect 8694 12315 8722 12334
rect 8750 12305 8778 12502
rect 8918 12417 8946 12423
rect 8918 12391 8919 12417
rect 8945 12391 8946 12417
rect 8750 12279 8751 12305
rect 8777 12279 8778 12305
rect 8750 12273 8778 12279
rect 8806 12361 8834 12367
rect 8806 12335 8807 12361
rect 8833 12335 8834 12361
rect 8358 11943 8359 11969
rect 8385 11943 8386 11969
rect 8358 11937 8386 11943
rect 8470 12138 8498 12143
rect 8470 11969 8498 12110
rect 8806 12138 8834 12335
rect 8806 12105 8834 12110
rect 8470 11943 8471 11969
rect 8497 11943 8498 11969
rect 8470 11937 8498 11943
rect 8918 11802 8946 12391
rect 8302 11718 8386 11746
rect 8078 11545 8106 11550
rect 8246 11577 8274 11583
rect 8246 11551 8247 11577
rect 8273 11551 8274 11577
rect 8134 11521 8162 11527
rect 8134 11495 8135 11521
rect 8161 11495 8162 11521
rect 8022 11465 8050 11471
rect 8022 11439 8023 11465
rect 8049 11439 8050 11465
rect 7574 11297 7658 11298
rect 7574 11271 7575 11297
rect 7601 11271 7658 11297
rect 7574 11270 7658 11271
rect 7966 11298 7994 11303
rect 8022 11298 8050 11439
rect 8134 11466 8162 11495
rect 8134 11433 8162 11438
rect 7966 11297 8050 11298
rect 7966 11271 7967 11297
rect 7993 11271 8050 11297
rect 7966 11270 8050 11271
rect 7574 11265 7602 11270
rect 7966 11265 7994 11270
rect 7490 11046 7546 11074
rect 7574 11130 7602 11135
rect 7462 11027 7490 11046
rect 7182 10794 7210 10799
rect 7182 10747 7210 10766
rect 7574 10794 7602 11102
rect 7910 11129 7938 11135
rect 7910 11103 7911 11129
rect 7937 11103 7938 11129
rect 6230 10738 6258 10743
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2086 10369 2114 10374
rect 6230 10401 6258 10710
rect 6846 10738 6874 10743
rect 6846 10691 6874 10710
rect 7294 10737 7322 10743
rect 7294 10711 7295 10737
rect 7321 10711 7322 10737
rect 6230 10375 6231 10401
rect 6257 10375 6258 10401
rect 6230 10369 6258 10375
rect 7070 10458 7098 10463
rect 7070 10345 7098 10430
rect 7238 10402 7266 10407
rect 7238 10355 7266 10374
rect 7070 10319 7071 10345
rect 7097 10319 7098 10345
rect 6062 10290 6090 10295
rect 5838 10289 6090 10290
rect 5838 10263 6063 10289
rect 6089 10263 6090 10289
rect 5838 10262 6090 10263
rect 5838 10065 5866 10262
rect 6062 10257 6090 10262
rect 5838 10039 5839 10065
rect 5865 10039 5866 10065
rect 5838 10033 5866 10039
rect 6006 10178 6034 10183
rect 5502 10010 5530 10015
rect 5502 10009 5642 10010
rect 5502 9983 5503 10009
rect 5529 9983 5642 10009
rect 5502 9982 5642 9983
rect 5502 9977 5530 9982
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 5614 9226 5642 9982
rect 5614 9179 5642 9198
rect 6006 9225 6034 10150
rect 7070 10178 7098 10319
rect 7294 10290 7322 10711
rect 7574 10737 7602 10766
rect 7574 10711 7575 10737
rect 7601 10711 7602 10737
rect 7574 10705 7602 10711
rect 7798 10793 7826 10799
rect 7798 10767 7799 10793
rect 7825 10767 7826 10793
rect 7518 10401 7546 10407
rect 7518 10375 7519 10401
rect 7545 10375 7546 10401
rect 7406 10290 7434 10295
rect 7294 10289 7434 10290
rect 7294 10263 7407 10289
rect 7433 10263 7434 10289
rect 7294 10262 7434 10263
rect 7070 10145 7098 10150
rect 7406 10122 7434 10262
rect 7406 10089 7434 10094
rect 7294 10010 7322 10015
rect 6902 10009 7378 10010
rect 6902 9983 7295 10009
rect 7321 9983 7378 10009
rect 6902 9982 7378 9983
rect 6902 9953 6930 9982
rect 7294 9977 7322 9982
rect 6902 9927 6903 9953
rect 6929 9927 6930 9953
rect 6902 9921 6930 9927
rect 7350 9617 7378 9982
rect 7518 9954 7546 10375
rect 7798 10402 7826 10767
rect 7910 10738 7938 11103
rect 8246 11130 8274 11551
rect 8246 11097 8274 11102
rect 7910 10705 7938 10710
rect 7966 11073 7994 11079
rect 7966 11047 7967 11073
rect 7993 11047 7994 11073
rect 7854 10402 7882 10407
rect 7798 10374 7854 10402
rect 7854 10065 7882 10374
rect 7854 10039 7855 10065
rect 7881 10039 7882 10065
rect 7518 9907 7546 9926
rect 7686 10009 7714 10015
rect 7686 9983 7687 10009
rect 7713 9983 7714 10009
rect 7350 9591 7351 9617
rect 7377 9591 7378 9617
rect 7350 9585 7378 9591
rect 7518 9562 7546 9567
rect 7518 9515 7546 9534
rect 7014 9505 7042 9511
rect 7014 9479 7015 9505
rect 7041 9479 7042 9505
rect 6006 9199 6007 9225
rect 6033 9199 6034 9225
rect 6006 9193 6034 9199
rect 6790 9226 6818 9231
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 6734 8442 6762 8447
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8073 994 8078
rect 6734 8106 6762 8414
rect 6790 8441 6818 9198
rect 7014 9226 7042 9479
rect 7014 9193 7042 9198
rect 7070 9506 7098 9511
rect 7070 9169 7098 9478
rect 7406 9506 7434 9511
rect 7406 9459 7434 9478
rect 7686 9506 7714 9983
rect 7854 9898 7882 10039
rect 7966 10010 7994 11047
rect 8190 10793 8218 10799
rect 8190 10767 8191 10793
rect 8217 10767 8218 10793
rect 8190 10738 8218 10767
rect 8190 10705 8218 10710
rect 8302 10793 8330 10799
rect 8302 10767 8303 10793
rect 8329 10767 8330 10793
rect 8302 10122 8330 10767
rect 8358 10737 8386 11718
rect 8526 11634 8554 11639
rect 8358 10711 8359 10737
rect 8385 10711 8386 10737
rect 8358 10705 8386 10711
rect 8414 10849 8442 10855
rect 8414 10823 8415 10849
rect 8441 10823 8442 10849
rect 8414 10290 8442 10823
rect 8302 10094 8386 10122
rect 8078 10066 8106 10071
rect 8078 10019 8106 10038
rect 7966 9977 7994 9982
rect 8302 10010 8330 10015
rect 8302 9963 8330 9982
rect 8022 9954 8050 9959
rect 8022 9907 8050 9926
rect 7854 9865 7882 9870
rect 8358 9730 8386 10094
rect 8358 9697 8386 9702
rect 8414 10065 8442 10262
rect 8414 10039 8415 10065
rect 8441 10039 8442 10065
rect 7686 9473 7714 9478
rect 8358 9617 8386 9623
rect 8358 9591 8359 9617
rect 8385 9591 8386 9617
rect 8358 9506 8386 9591
rect 8358 9473 8386 9478
rect 8414 9338 8442 10039
rect 8526 10457 8554 11606
rect 8918 11578 8946 11774
rect 9366 11689 9394 12614
rect 9534 12025 9562 13119
rect 9926 13145 9954 13151
rect 9926 13119 9927 13145
rect 9953 13119 9954 13145
rect 9926 12698 9954 13119
rect 9814 12670 9954 12698
rect 10542 13145 10570 13151
rect 10542 13119 10543 13145
rect 10569 13119 10570 13145
rect 9814 12474 9842 12670
rect 10542 12586 10570 13119
rect 10766 12809 10794 13399
rect 10878 13201 10906 13566
rect 10878 13175 10879 13201
rect 10905 13175 10906 13201
rect 10878 13169 10906 13175
rect 10766 12783 10767 12809
rect 10793 12783 10794 12809
rect 10766 12777 10794 12783
rect 11942 13089 11970 15946
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 18830 13538 18858 13543
rect 18774 13537 18858 13538
rect 18774 13511 18831 13537
rect 18857 13511 18858 13537
rect 18774 13510 18858 13511
rect 13062 13201 13090 13207
rect 13062 13175 13063 13201
rect 13089 13175 13090 13201
rect 12838 13145 12866 13151
rect 12838 13119 12839 13145
rect 12865 13119 12866 13145
rect 11942 13063 11943 13089
rect 11969 13063 11970 13089
rect 10990 12754 11018 12759
rect 10990 12707 11018 12726
rect 11942 12754 11970 13063
rect 12222 13089 12250 13095
rect 12222 13063 12223 13089
rect 12249 13063 12250 13089
rect 11942 12721 11970 12726
rect 12110 12754 12138 12759
rect 12222 12754 12250 13063
rect 12110 12753 12250 12754
rect 12110 12727 12111 12753
rect 12137 12727 12250 12753
rect 12110 12726 12250 12727
rect 12110 12721 12138 12726
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10542 12553 10570 12558
rect 10710 12641 10738 12647
rect 10710 12615 10711 12641
rect 10737 12615 10738 12641
rect 9918 12525 10050 12530
rect 9870 12474 9898 12479
rect 9814 12473 9898 12474
rect 9814 12447 9871 12473
rect 9897 12447 9898 12473
rect 9814 12446 9898 12447
rect 9870 12441 9898 12446
rect 9926 12417 9954 12423
rect 9926 12391 9927 12417
rect 9953 12391 9954 12417
rect 9534 11999 9535 12025
rect 9561 11999 9562 12025
rect 9534 11993 9562 11999
rect 9814 12362 9842 12367
rect 9590 11970 9618 11975
rect 9478 11914 9506 11933
rect 9478 11881 9506 11886
rect 9534 11913 9562 11919
rect 9534 11887 9535 11913
rect 9561 11887 9562 11913
rect 9478 11802 9506 11807
rect 9534 11802 9562 11887
rect 9590 11913 9618 11942
rect 9590 11887 9591 11913
rect 9617 11887 9618 11913
rect 9590 11881 9618 11887
rect 9814 11914 9842 12334
rect 9926 12138 9954 12391
rect 9926 12105 9954 12110
rect 10038 12361 10066 12367
rect 10038 12335 10039 12361
rect 10065 12335 10066 12361
rect 9506 11774 9562 11802
rect 9702 11857 9730 11863
rect 9702 11831 9703 11857
rect 9729 11831 9730 11857
rect 9478 11769 9506 11774
rect 9366 11663 9367 11689
rect 9393 11663 9394 11689
rect 9366 11657 9394 11663
rect 9702 11690 9730 11831
rect 9702 11657 9730 11662
rect 9142 11634 9170 11639
rect 9086 11633 9170 11634
rect 9086 11607 9143 11633
rect 9169 11607 9170 11633
rect 9086 11606 9170 11607
rect 9030 11578 9058 11583
rect 8918 11577 9058 11578
rect 8918 11551 9031 11577
rect 9057 11551 9058 11577
rect 8918 11550 9058 11551
rect 8750 11466 8778 11471
rect 8526 10431 8527 10457
rect 8553 10431 8554 10457
rect 8470 9505 8498 9511
rect 8470 9479 8471 9505
rect 8497 9479 8498 9505
rect 8470 9450 8498 9479
rect 8470 9417 8498 9422
rect 8414 9305 8442 9310
rect 7294 9226 7322 9231
rect 8526 9226 8554 10431
rect 8694 11438 8750 11466
rect 8638 10010 8666 10015
rect 8638 9963 8666 9982
rect 7294 9179 7322 9198
rect 8414 9198 8526 9226
rect 7070 9143 7071 9169
rect 7097 9143 7098 9169
rect 7070 9137 7098 9143
rect 8190 8834 8218 8839
rect 7126 8722 7154 8727
rect 7126 8497 7154 8694
rect 7126 8471 7127 8497
rect 7153 8471 7154 8497
rect 7126 8465 7154 8471
rect 7798 8554 7826 8559
rect 6790 8415 6791 8441
rect 6817 8415 6818 8441
rect 6790 8409 6818 8415
rect 6734 8059 6762 8078
rect 7798 8105 7826 8526
rect 8190 8385 8218 8806
rect 8358 8722 8386 8727
rect 8358 8675 8386 8694
rect 8414 8554 8442 9198
rect 8526 9193 8554 9198
rect 8582 9730 8610 9735
rect 8694 9730 8722 11438
rect 8750 11433 8778 11438
rect 8918 10794 8946 10799
rect 8918 10793 9002 10794
rect 8918 10767 8919 10793
rect 8945 10767 9002 10793
rect 8918 10766 9002 10767
rect 8918 10761 8946 10766
rect 8806 10066 8834 10071
rect 8974 10066 9002 10766
rect 8806 10065 8890 10066
rect 8806 10039 8807 10065
rect 8833 10039 8890 10065
rect 8806 10038 8890 10039
rect 8806 10033 8834 10038
rect 8526 8834 8554 8839
rect 8582 8834 8610 9702
rect 8638 9702 8722 9730
rect 8750 10009 8778 10015
rect 8750 9983 8751 10009
rect 8777 9983 8778 10009
rect 8638 9170 8666 9702
rect 8750 9674 8778 9983
rect 8862 9786 8890 10038
rect 8974 10009 9002 10038
rect 8974 9983 8975 10009
rect 9001 9983 9002 10009
rect 8974 9977 9002 9983
rect 9030 9898 9058 11550
rect 8862 9753 8890 9758
rect 8918 9870 9058 9898
rect 8750 9646 8834 9674
rect 8694 9618 8722 9623
rect 8806 9618 8834 9646
rect 8694 9617 8778 9618
rect 8694 9591 8695 9617
rect 8721 9591 8778 9617
rect 8694 9590 8778 9591
rect 8806 9590 8890 9618
rect 8694 9585 8722 9590
rect 8750 9282 8778 9590
rect 8806 9505 8834 9511
rect 8806 9479 8807 9505
rect 8833 9479 8834 9505
rect 8806 9338 8834 9479
rect 8806 9305 8834 9310
rect 8750 9235 8778 9254
rect 8638 9137 8666 9142
rect 8694 9226 8722 9231
rect 8694 9058 8722 9198
rect 8526 8833 8610 8834
rect 8526 8807 8527 8833
rect 8553 8807 8610 8833
rect 8526 8806 8610 8807
rect 8638 9030 8722 9058
rect 8806 9169 8834 9175
rect 8806 9143 8807 9169
rect 8833 9143 8834 9169
rect 8638 8890 8666 9030
rect 8470 8722 8498 8727
rect 8470 8675 8498 8694
rect 8526 8610 8554 8806
rect 8190 8359 8191 8385
rect 8217 8359 8218 8385
rect 8190 8353 8218 8359
rect 8246 8553 8442 8554
rect 8246 8527 8415 8553
rect 8441 8527 8442 8553
rect 8246 8526 8442 8527
rect 7798 8079 7799 8105
rect 7825 8079 7826 8105
rect 7798 8073 7826 8079
rect 8190 8050 8218 8055
rect 8246 8050 8274 8526
rect 8414 8521 8442 8526
rect 8470 8582 8554 8610
rect 8190 8049 8274 8050
rect 8190 8023 8191 8049
rect 8217 8023 8274 8049
rect 8190 8022 8274 8023
rect 8190 8017 8218 8022
rect 8246 7770 8274 8022
rect 8358 8050 8386 8055
rect 8358 8003 8386 8022
rect 8302 7770 8330 7775
rect 8246 7769 8330 7770
rect 8246 7743 8303 7769
rect 8329 7743 8330 7769
rect 8246 7742 8330 7743
rect 8134 7602 8162 7607
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 8134 7321 8162 7574
rect 8134 7295 8135 7321
rect 8161 7295 8162 7321
rect 8134 7289 8162 7295
rect 7798 7266 7826 7271
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 7798 6481 7826 7238
rect 8246 7266 8274 7742
rect 8302 7737 8330 7742
rect 8246 7233 8274 7238
rect 8470 7210 8498 8582
rect 8526 8106 8554 8111
rect 8526 8049 8554 8078
rect 8526 8023 8527 8049
rect 8553 8023 8554 8049
rect 8526 8017 8554 8023
rect 8638 8049 8666 8862
rect 8750 8834 8778 8839
rect 8806 8834 8834 9143
rect 8778 8806 8834 8834
rect 8750 8787 8778 8806
rect 8862 8778 8890 9590
rect 8862 8731 8890 8750
rect 8694 8554 8722 8559
rect 8694 8507 8722 8526
rect 8806 8498 8834 8503
rect 8806 8442 8834 8470
rect 8806 8441 8890 8442
rect 8806 8415 8807 8441
rect 8833 8415 8890 8441
rect 8806 8414 8890 8415
rect 8806 8409 8834 8414
rect 8806 8330 8834 8335
rect 8638 8023 8639 8049
rect 8665 8023 8666 8049
rect 8638 8017 8666 8023
rect 8694 8329 8834 8330
rect 8694 8303 8807 8329
rect 8833 8303 8834 8329
rect 8694 8302 8834 8303
rect 8582 7938 8610 7943
rect 8694 7938 8722 8302
rect 8806 8297 8834 8302
rect 8862 8162 8890 8414
rect 8582 7937 8722 7938
rect 8582 7911 8583 7937
rect 8609 7911 8722 7937
rect 8582 7910 8722 7911
rect 8806 8134 8890 8162
rect 8582 7905 8610 7910
rect 8806 7657 8834 8134
rect 8806 7631 8807 7657
rect 8833 7631 8834 7657
rect 8806 7625 8834 7631
rect 8918 7657 8946 9870
rect 9086 9730 9114 11606
rect 9142 11601 9170 11606
rect 9198 11634 9226 11639
rect 9198 11587 9226 11606
rect 9758 11634 9786 11639
rect 9534 11577 9562 11583
rect 9534 11551 9535 11577
rect 9561 11551 9562 11577
rect 9142 11186 9170 11191
rect 9142 10849 9170 11158
rect 9478 11185 9506 11191
rect 9478 11159 9479 11185
rect 9505 11159 9506 11185
rect 9366 11074 9394 11079
rect 9366 11027 9394 11046
rect 9142 10823 9143 10849
rect 9169 10823 9170 10849
rect 9142 10817 9170 10823
rect 9478 10570 9506 11159
rect 9478 10537 9506 10542
rect 9534 10794 9562 11551
rect 9702 11578 9730 11583
rect 9590 11186 9618 11191
rect 9702 11186 9730 11550
rect 9618 11158 9730 11186
rect 9590 11139 9618 11158
rect 9758 10849 9786 11606
rect 9814 10905 9842 11886
rect 10038 11858 10066 12335
rect 10150 12362 10178 12367
rect 10150 12315 10178 12334
rect 10542 12138 10570 12143
rect 10094 11970 10122 11975
rect 10094 11969 10346 11970
rect 10094 11943 10095 11969
rect 10121 11943 10346 11969
rect 10094 11942 10346 11943
rect 10094 11937 10122 11942
rect 10150 11858 10178 11863
rect 10038 11825 10066 11830
rect 10094 11857 10178 11858
rect 10094 11831 10151 11857
rect 10177 11831 10178 11857
rect 10094 11830 10178 11831
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9870 11690 9898 11695
rect 9870 11129 9898 11662
rect 10094 11634 10122 11830
rect 10150 11825 10178 11830
rect 10262 11858 10290 11863
rect 10262 11811 10290 11830
rect 10094 11587 10122 11606
rect 9926 11577 9954 11583
rect 9926 11551 9927 11577
rect 9953 11551 9954 11577
rect 9926 11522 9954 11551
rect 9926 11489 9954 11494
rect 10318 11466 10346 11942
rect 10542 11689 10570 12110
rect 10542 11663 10543 11689
rect 10569 11663 10570 11689
rect 10542 11657 10570 11663
rect 10318 11186 10346 11438
rect 10318 11153 10346 11158
rect 10374 11633 10402 11639
rect 10374 11607 10375 11633
rect 10401 11607 10402 11633
rect 10374 11522 10402 11607
rect 10654 11633 10682 11639
rect 10654 11607 10655 11633
rect 10681 11607 10682 11633
rect 10654 11578 10682 11607
rect 10710 11634 10738 12615
rect 10766 12641 10794 12647
rect 10766 12615 10767 12641
rect 10793 12615 10794 12641
rect 10766 11970 10794 12615
rect 10878 12642 10906 12647
rect 10878 12595 10906 12614
rect 10766 11937 10794 11942
rect 11270 12586 11298 12591
rect 11270 11969 11298 12558
rect 12222 12586 12250 12726
rect 12222 12553 12250 12558
rect 12446 12697 12474 12703
rect 12446 12671 12447 12697
rect 12473 12671 12474 12697
rect 12446 12082 12474 12671
rect 12782 12586 12810 12591
rect 12782 12473 12810 12558
rect 12782 12447 12783 12473
rect 12809 12447 12810 12473
rect 12782 12418 12810 12447
rect 12782 12385 12810 12390
rect 12838 12250 12866 13119
rect 12950 13146 12978 13151
rect 12950 13145 13034 13146
rect 12950 13119 12951 13145
rect 12977 13119 13034 13145
rect 12950 13118 13034 13119
rect 12950 13113 12978 13118
rect 12894 13034 12922 13039
rect 12894 13033 12978 13034
rect 12894 13007 12895 13033
rect 12921 13007 12978 13033
rect 12894 13006 12978 13007
rect 12894 13001 12922 13006
rect 12838 12217 12866 12222
rect 12446 12049 12474 12054
rect 12782 12082 12810 12087
rect 12670 12026 12698 12031
rect 11270 11943 11271 11969
rect 11297 11943 11298 11969
rect 11270 11937 11298 11943
rect 11550 11970 11578 11975
rect 11550 11802 11578 11942
rect 11606 11914 11634 11919
rect 11606 11913 11746 11914
rect 11606 11887 11607 11913
rect 11633 11887 11746 11913
rect 11606 11886 11746 11887
rect 11606 11881 11634 11886
rect 11550 11774 11634 11802
rect 10934 11746 10962 11751
rect 10710 11606 10850 11634
rect 10822 11578 10850 11606
rect 10682 11550 10794 11578
rect 10654 11545 10682 11550
rect 9870 11103 9871 11129
rect 9897 11103 9898 11129
rect 9870 11074 9898 11103
rect 9870 11046 10122 11074
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9814 10879 9815 10905
rect 9841 10879 9842 10905
rect 9814 10873 9842 10879
rect 9758 10823 9759 10849
rect 9785 10823 9786 10849
rect 9758 10817 9786 10823
rect 9310 10010 9338 10015
rect 8974 9702 9114 9730
rect 9198 10009 9338 10010
rect 9198 9983 9311 10009
rect 9337 9983 9338 10009
rect 9198 9982 9338 9983
rect 9198 9898 9226 9982
rect 9310 9977 9338 9982
rect 8974 9282 9002 9702
rect 9030 9618 9058 9623
rect 9198 9618 9226 9870
rect 9030 9617 9226 9618
rect 9030 9591 9031 9617
rect 9057 9591 9226 9617
rect 9030 9590 9226 9591
rect 9254 9617 9282 9623
rect 9254 9591 9255 9617
rect 9281 9591 9282 9617
rect 9030 9585 9058 9590
rect 9254 9562 9282 9591
rect 9254 9529 9282 9534
rect 9478 9506 9506 9511
rect 9142 9450 9170 9455
rect 8974 9254 9058 9282
rect 8974 9170 9002 9175
rect 8974 8834 9002 9142
rect 9030 8946 9058 9254
rect 9030 8913 9058 8918
rect 9086 9114 9114 9119
rect 8974 8806 9058 8834
rect 8974 8722 9002 8727
rect 8974 8554 9002 8694
rect 9030 8666 9058 8806
rect 9086 8778 9114 9086
rect 9142 8833 9170 9422
rect 9254 9226 9282 9231
rect 9254 9179 9282 9198
rect 9422 9226 9450 9231
rect 9422 8889 9450 9198
rect 9478 9225 9506 9478
rect 9534 9450 9562 10766
rect 9814 10793 9842 10799
rect 9814 10767 9815 10793
rect 9841 10767 9842 10793
rect 9702 10010 9730 10015
rect 9590 10009 9730 10010
rect 9590 9983 9703 10009
rect 9729 9983 9730 10009
rect 9590 9982 9730 9983
rect 9590 9954 9618 9982
rect 9702 9977 9730 9982
rect 9590 9561 9618 9926
rect 9590 9535 9591 9561
rect 9617 9535 9618 9561
rect 9590 9529 9618 9535
rect 9702 9730 9730 9735
rect 9702 9505 9730 9702
rect 9702 9479 9703 9505
rect 9729 9479 9730 9505
rect 9702 9473 9730 9479
rect 9814 9674 9842 10767
rect 10094 10682 10122 11046
rect 10094 10649 10122 10654
rect 10038 10401 10066 10407
rect 10038 10375 10039 10401
rect 10065 10375 10066 10401
rect 10038 10346 10066 10375
rect 10038 10313 10066 10318
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10206 10066 10234 10071
rect 10206 9730 10234 10038
rect 10206 9683 10234 9702
rect 9814 9646 9954 9674
rect 9534 9422 9618 9450
rect 9534 9282 9562 9287
rect 9534 9235 9562 9254
rect 9478 9199 9479 9225
rect 9505 9199 9506 9225
rect 9478 9193 9506 9199
rect 9590 9169 9618 9422
rect 9814 9226 9842 9646
rect 9926 9617 9954 9646
rect 9926 9591 9927 9617
rect 9953 9591 9954 9617
rect 9926 9585 9954 9591
rect 10318 9673 10346 9679
rect 10318 9647 10319 9673
rect 10345 9647 10346 9673
rect 9870 9562 9898 9567
rect 9870 9515 9898 9534
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10262 9338 10290 9343
rect 10150 9282 10178 9287
rect 10094 9254 10150 9282
rect 10038 9226 10066 9231
rect 9814 9193 9842 9198
rect 9982 9198 10038 9226
rect 9590 9143 9591 9169
rect 9617 9143 9618 9169
rect 9590 9137 9618 9143
rect 9982 8945 10010 9198
rect 10038 9179 10066 9198
rect 10094 9114 10122 9254
rect 10150 9249 10178 9254
rect 10262 9226 10290 9310
rect 9982 8919 9983 8945
rect 10009 8919 10010 8945
rect 9982 8913 10010 8919
rect 10038 9086 10122 9114
rect 10206 9225 10290 9226
rect 10206 9199 10263 9225
rect 10289 9199 10290 9225
rect 10206 9198 10290 9199
rect 9422 8863 9423 8889
rect 9449 8863 9450 8889
rect 9422 8857 9450 8863
rect 10038 8889 10066 9086
rect 10206 8945 10234 9198
rect 10262 9193 10290 9198
rect 10206 8919 10207 8945
rect 10233 8919 10234 8945
rect 10206 8913 10234 8919
rect 10262 8946 10290 8951
rect 10038 8863 10039 8889
rect 10065 8863 10066 8889
rect 9142 8807 9143 8833
rect 9169 8807 9170 8833
rect 9142 8801 9170 8807
rect 9478 8834 9506 8839
rect 9478 8787 9506 8806
rect 9702 8834 9730 8839
rect 10038 8834 10066 8863
rect 10262 8889 10290 8918
rect 10262 8863 10263 8889
rect 10289 8863 10290 8889
rect 10262 8857 10290 8863
rect 9702 8833 10066 8834
rect 9702 8807 9703 8833
rect 9729 8807 10066 8833
rect 9702 8806 10066 8807
rect 9702 8801 9730 8806
rect 9086 8731 9114 8750
rect 10318 8778 10346 9647
rect 10374 9617 10402 11494
rect 10654 11186 10682 11191
rect 10654 11139 10682 11158
rect 10766 11129 10794 11550
rect 10822 11531 10850 11550
rect 10766 11103 10767 11129
rect 10793 11103 10794 11129
rect 10766 11097 10794 11103
rect 10934 11186 10962 11718
rect 10934 11073 10962 11158
rect 11326 11578 11354 11583
rect 11102 11130 11130 11135
rect 11102 11083 11130 11102
rect 10934 11047 10935 11073
rect 10961 11047 10962 11073
rect 10934 11041 10962 11047
rect 10486 10794 10514 10799
rect 10486 10747 10514 10766
rect 11158 10793 11186 10799
rect 11158 10767 11159 10793
rect 11185 10767 11186 10793
rect 10766 10738 10794 10743
rect 10430 10682 10458 10687
rect 10458 10654 10514 10682
rect 10430 10649 10458 10654
rect 10430 10570 10458 10575
rect 10430 10065 10458 10542
rect 10430 10039 10431 10065
rect 10457 10039 10458 10065
rect 10430 10033 10458 10039
rect 10374 9591 10375 9617
rect 10401 9591 10402 9617
rect 10374 9562 10402 9591
rect 10374 9529 10402 9534
rect 10374 9170 10402 9175
rect 10486 9170 10514 10654
rect 10542 10066 10570 10071
rect 10542 9282 10570 10038
rect 10766 9953 10794 10710
rect 10934 10402 10962 10407
rect 10934 10355 10962 10374
rect 11046 10065 11074 10071
rect 11046 10039 11047 10065
rect 11073 10039 11074 10065
rect 10766 9927 10767 9953
rect 10793 9927 10794 9953
rect 10766 9921 10794 9927
rect 10934 10009 10962 10015
rect 10934 9983 10935 10009
rect 10961 9983 10962 10009
rect 10934 9617 10962 9983
rect 10934 9591 10935 9617
rect 10961 9591 10962 9617
rect 10934 9282 10962 9591
rect 10990 9673 11018 9679
rect 10990 9647 10991 9673
rect 11017 9647 11018 9673
rect 10990 9618 11018 9647
rect 10990 9585 11018 9590
rect 10542 9235 10570 9254
rect 10878 9254 10962 9282
rect 10374 8833 10402 9142
rect 10374 8807 10375 8833
rect 10401 8807 10402 8833
rect 10374 8801 10402 8807
rect 10430 9169 10514 9170
rect 10430 9143 10487 9169
rect 10513 9143 10514 9169
rect 10430 9142 10514 9143
rect 9030 8638 9114 8666
rect 8974 8526 9058 8554
rect 8974 8441 9002 8447
rect 8974 8415 8975 8441
rect 9001 8415 9002 8441
rect 8974 8386 9002 8415
rect 9030 8442 9058 8526
rect 9086 8497 9114 8638
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9086 8471 9087 8497
rect 9113 8471 9114 8497
rect 9086 8465 9114 8471
rect 9254 8498 9282 8503
rect 9254 8451 9282 8470
rect 9030 8409 9058 8414
rect 9534 8442 9562 8447
rect 9534 8395 9562 8414
rect 8974 8353 9002 8358
rect 8918 7631 8919 7657
rect 8945 7631 8946 7657
rect 8918 7625 8946 7631
rect 9030 8330 9058 8335
rect 8974 7602 9002 7621
rect 8974 7569 9002 7574
rect 8470 7177 8498 7182
rect 8974 7210 9002 7215
rect 8806 6930 8834 6935
rect 8806 6929 8946 6930
rect 8806 6903 8807 6929
rect 8833 6903 8946 6929
rect 8806 6902 8946 6903
rect 8806 6897 8834 6902
rect 8134 6818 8162 6823
rect 8134 6537 8162 6790
rect 8862 6818 8890 6823
rect 8862 6771 8890 6790
rect 8918 6762 8946 6902
rect 8974 6929 9002 7182
rect 8974 6903 8975 6929
rect 9001 6903 9002 6929
rect 8974 6897 9002 6903
rect 9030 6873 9058 8302
rect 9422 8330 9450 8335
rect 9422 8283 9450 8302
rect 10318 8162 10346 8750
rect 10374 8162 10402 8167
rect 10318 8161 10402 8162
rect 10318 8135 10375 8161
rect 10401 8135 10402 8161
rect 10318 8134 10402 8135
rect 10374 8129 10402 8134
rect 10430 8050 10458 9142
rect 10486 9137 10514 9142
rect 10766 9226 10794 9231
rect 10766 8834 10794 9198
rect 10766 8801 10794 8806
rect 10822 9169 10850 9175
rect 10822 9143 10823 9169
rect 10849 9143 10850 9169
rect 10822 8945 10850 9143
rect 10878 9170 10906 9254
rect 10990 9226 11018 9231
rect 10878 9137 10906 9142
rect 10934 9170 10962 9175
rect 10990 9170 11018 9198
rect 10934 9169 11018 9170
rect 10934 9143 10935 9169
rect 10961 9143 11018 9169
rect 10934 9142 11018 9143
rect 10934 9114 10962 9142
rect 11046 9114 11074 10039
rect 11158 9729 11186 10767
rect 11158 9703 11159 9729
rect 11185 9703 11186 9729
rect 11158 9697 11186 9703
rect 11102 9617 11130 9623
rect 11102 9591 11103 9617
rect 11129 9591 11130 9617
rect 11102 9338 11130 9591
rect 11102 9291 11130 9310
rect 11326 9282 11354 11550
rect 11550 11578 11578 11583
rect 11550 11531 11578 11550
rect 11382 11241 11410 11247
rect 11382 11215 11383 11241
rect 11409 11215 11410 11241
rect 11382 10066 11410 11215
rect 11606 10849 11634 11774
rect 11718 11690 11746 11886
rect 11774 11690 11802 11695
rect 11718 11689 11802 11690
rect 11718 11663 11775 11689
rect 11801 11663 11802 11689
rect 11718 11662 11802 11663
rect 11774 11657 11802 11662
rect 12670 11689 12698 11998
rect 12782 11969 12810 12054
rect 12782 11943 12783 11969
rect 12809 11943 12810 11969
rect 12782 11937 12810 11943
rect 12950 11969 12978 13006
rect 13006 12530 13034 13118
rect 13062 12810 13090 13175
rect 13678 13089 13706 13095
rect 13678 13063 13679 13089
rect 13705 13063 13706 13089
rect 13062 12777 13090 12782
rect 13510 12810 13538 12815
rect 13510 12763 13538 12782
rect 13342 12698 13370 12703
rect 13006 12502 13314 12530
rect 12950 11943 12951 11969
rect 12977 11943 12978 11969
rect 12950 11937 12978 11943
rect 13006 12418 13034 12423
rect 13006 12361 13034 12390
rect 13006 12335 13007 12361
rect 13033 12335 13034 12361
rect 12894 11858 12922 11863
rect 12894 11811 12922 11830
rect 12782 11802 12810 11807
rect 12670 11663 12671 11689
rect 12697 11663 12698 11689
rect 12670 11657 12698 11663
rect 12726 11774 12782 11802
rect 12726 11633 12754 11774
rect 12782 11769 12810 11774
rect 12950 11690 12978 11695
rect 13006 11690 13034 12335
rect 13118 12250 13146 12255
rect 13146 12222 13202 12250
rect 13118 12217 13146 12222
rect 12726 11607 12727 11633
rect 12753 11607 12754 11633
rect 11718 11577 11746 11583
rect 11718 11551 11719 11577
rect 11745 11551 11746 11577
rect 11718 10906 11746 11551
rect 11886 11578 11914 11583
rect 11886 11531 11914 11550
rect 12558 11578 12586 11583
rect 12558 11531 12586 11550
rect 12726 11354 12754 11607
rect 12614 11326 12754 11354
rect 12838 11689 13034 11690
rect 12838 11663 12951 11689
rect 12977 11663 13034 11689
rect 12838 11662 13034 11663
rect 13174 11969 13202 12222
rect 13174 11943 13175 11969
rect 13201 11943 13202 11969
rect 11886 11130 11914 11135
rect 12446 11130 12474 11135
rect 11718 10878 11858 10906
rect 11606 10823 11607 10849
rect 11633 10823 11634 10849
rect 11550 10402 11578 10407
rect 11550 10121 11578 10374
rect 11550 10095 11551 10121
rect 11577 10095 11578 10121
rect 11550 10089 11578 10095
rect 11382 10033 11410 10038
rect 11326 9254 11410 9282
rect 11326 9169 11354 9175
rect 11326 9143 11327 9169
rect 11353 9143 11354 9169
rect 11326 9114 11354 9143
rect 11046 9086 11354 9114
rect 10934 9081 10962 9086
rect 10822 8919 10823 8945
rect 10849 8919 10850 8945
rect 10654 8721 10682 8727
rect 10654 8695 10655 8721
rect 10681 8695 10682 8721
rect 10654 8610 10682 8695
rect 10598 8582 10654 8610
rect 10598 8330 10626 8582
rect 10654 8577 10682 8582
rect 10822 8553 10850 8919
rect 10934 8946 10962 8951
rect 10934 8889 10962 8918
rect 10934 8863 10935 8889
rect 10961 8863 10962 8889
rect 10934 8857 10962 8863
rect 11102 8834 11130 8839
rect 11102 8787 11130 8806
rect 10822 8527 10823 8553
rect 10849 8527 10850 8553
rect 10822 8521 10850 8527
rect 10654 8497 10682 8503
rect 10654 8471 10655 8497
rect 10681 8471 10682 8497
rect 10654 8386 10682 8471
rect 10654 8353 10682 8358
rect 10598 8297 10626 8302
rect 11158 8330 11186 9086
rect 11382 9002 11410 9254
rect 11214 8974 11410 9002
rect 11494 9225 11522 9231
rect 11494 9199 11495 9225
rect 11521 9199 11522 9225
rect 11214 8497 11242 8974
rect 11494 8946 11522 9199
rect 11494 8913 11522 8918
rect 11382 8890 11410 8895
rect 11382 8843 11410 8862
rect 11214 8471 11215 8497
rect 11241 8471 11242 8497
rect 11214 8386 11242 8471
rect 11382 8442 11410 8447
rect 11382 8395 11410 8414
rect 11494 8441 11522 8447
rect 11494 8415 11495 8441
rect 11521 8415 11522 8441
rect 11214 8353 11242 8358
rect 11270 8385 11298 8391
rect 11270 8359 11271 8385
rect 11297 8359 11298 8385
rect 11158 8297 11186 8302
rect 11270 8105 11298 8359
rect 11270 8079 11271 8105
rect 11297 8079 11298 8105
rect 11270 8073 11298 8079
rect 11494 8106 11522 8415
rect 11606 8442 11634 10823
rect 11830 10850 11858 10878
rect 11774 10794 11802 10799
rect 11662 10793 11802 10794
rect 11662 10767 11775 10793
rect 11801 10767 11802 10793
rect 11662 10766 11802 10767
rect 11662 9730 11690 10766
rect 11774 10761 11802 10766
rect 11830 10682 11858 10822
rect 11662 9337 11690 9702
rect 11662 9311 11663 9337
rect 11689 9311 11690 9337
rect 11662 9305 11690 9311
rect 11718 10654 11858 10682
rect 11718 9169 11746 10654
rect 11830 10346 11858 10351
rect 11774 10066 11802 10071
rect 11774 10019 11802 10038
rect 11830 9617 11858 10318
rect 11830 9591 11831 9617
rect 11857 9591 11858 9617
rect 11830 9585 11858 9591
rect 11774 9338 11802 9343
rect 11886 9338 11914 11102
rect 11942 11129 12474 11130
rect 11942 11103 12447 11129
rect 12473 11103 12474 11129
rect 11942 11102 12474 11103
rect 11942 10682 11970 11102
rect 12446 11097 12474 11102
rect 11998 10850 12026 10855
rect 11998 10803 12026 10822
rect 12054 10794 12082 10799
rect 12054 10793 12194 10794
rect 12054 10767 12055 10793
rect 12081 10767 12194 10793
rect 12054 10766 12194 10767
rect 12054 10761 12082 10766
rect 11998 10682 12026 10687
rect 11942 10681 12026 10682
rect 11942 10655 11999 10681
rect 12025 10655 12026 10681
rect 11942 10654 12026 10655
rect 11998 10649 12026 10654
rect 12166 10121 12194 10766
rect 12166 10095 12167 10121
rect 12193 10095 12194 10121
rect 12166 10089 12194 10095
rect 12278 10066 12306 10071
rect 12278 10019 12306 10038
rect 12614 10066 12642 11326
rect 12838 11185 12866 11662
rect 12950 11657 12978 11662
rect 13174 11354 13202 11943
rect 13286 11969 13314 12502
rect 13342 12025 13370 12670
rect 13622 12642 13650 12647
rect 13398 12641 13650 12642
rect 13398 12615 13623 12641
rect 13649 12615 13650 12641
rect 13398 12614 13650 12615
rect 13398 12417 13426 12614
rect 13622 12609 13650 12614
rect 13678 12586 13706 13063
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 14182 12753 14210 12759
rect 14182 12727 14183 12753
rect 14209 12727 14210 12753
rect 13790 12698 13818 12703
rect 13790 12651 13818 12670
rect 13678 12553 13706 12558
rect 13734 12641 13762 12647
rect 13734 12615 13735 12641
rect 13761 12615 13762 12641
rect 13398 12391 13399 12417
rect 13425 12391 13426 12417
rect 13398 12385 13426 12391
rect 13342 11999 13343 12025
rect 13369 11999 13370 12025
rect 13342 11993 13370 11999
rect 13398 12306 13426 12311
rect 13286 11943 13287 11969
rect 13313 11943 13314 11969
rect 13286 11802 13314 11943
rect 13398 11913 13426 12278
rect 13734 12138 13762 12615
rect 14182 12642 14210 12727
rect 14294 12698 14322 12703
rect 14294 12651 14322 12670
rect 14182 12609 14210 12614
rect 14574 12642 14602 12647
rect 14518 12306 14546 12311
rect 14574 12306 14602 12614
rect 14742 12642 14770 12647
rect 14742 12595 14770 12614
rect 18774 12642 18802 13510
rect 18830 13505 18858 13510
rect 18942 13145 18970 13151
rect 18942 13119 18943 13145
rect 18969 13119 18970 13145
rect 18830 12754 18858 12759
rect 18830 12707 18858 12726
rect 18942 12698 18970 13119
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 19950 13089 19978 13095
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 19950 12810 19978 13063
rect 19950 12777 19978 12782
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 18942 12665 18970 12670
rect 18774 12609 18802 12614
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 18830 12362 18858 12367
rect 18830 12315 18858 12334
rect 14546 12278 14602 12306
rect 14798 12305 14826 12311
rect 14798 12279 14799 12305
rect 14825 12279 14826 12305
rect 14518 12259 14546 12278
rect 13734 12105 13762 12110
rect 13398 11887 13399 11913
rect 13425 11887 13426 11913
rect 13398 11881 13426 11887
rect 13286 11769 13314 11774
rect 13174 11326 13426 11354
rect 13062 11298 13090 11303
rect 13062 11297 13202 11298
rect 13062 11271 13063 11297
rect 13089 11271 13202 11297
rect 13062 11270 13202 11271
rect 13062 11265 13090 11270
rect 12838 11159 12839 11185
rect 12865 11159 12866 11185
rect 12838 10906 12866 11159
rect 13118 11186 13146 11191
rect 13118 11139 13146 11158
rect 13006 11130 13034 11135
rect 12838 10793 12866 10878
rect 12838 10767 12839 10793
rect 12865 10767 12866 10793
rect 12838 10761 12866 10767
rect 12894 11129 13034 11130
rect 12894 11103 13007 11129
rect 13033 11103 13034 11129
rect 12894 11102 13034 11103
rect 12614 10019 12642 10038
rect 12894 10290 12922 11102
rect 13006 11097 13034 11102
rect 13174 10850 13202 11270
rect 13230 11270 13370 11298
rect 13230 11185 13258 11270
rect 13230 11159 13231 11185
rect 13257 11159 13258 11185
rect 13230 11153 13258 11159
rect 13286 11185 13314 11191
rect 13286 11159 13287 11185
rect 13313 11159 13314 11185
rect 13230 10850 13258 10855
rect 13174 10849 13258 10850
rect 13174 10823 13231 10849
rect 13257 10823 13258 10849
rect 13174 10822 13258 10823
rect 13230 10817 13258 10822
rect 12334 10009 12362 10015
rect 12334 9983 12335 10009
rect 12361 9983 12362 10009
rect 11998 9954 12026 9959
rect 11774 9337 11914 9338
rect 11774 9311 11775 9337
rect 11801 9311 11914 9337
rect 11774 9310 11914 9311
rect 11942 9953 12026 9954
rect 11942 9927 11999 9953
rect 12025 9927 12026 9953
rect 11942 9926 12026 9927
rect 11774 9305 11802 9310
rect 11718 9143 11719 9169
rect 11745 9143 11746 9169
rect 11718 9137 11746 9143
rect 11942 9225 11970 9926
rect 11998 9921 12026 9926
rect 12334 9618 12362 9983
rect 11942 9199 11943 9225
rect 11969 9199 11970 9225
rect 11942 9170 11970 9199
rect 11942 9137 11970 9142
rect 12110 9281 12138 9287
rect 12110 9255 12111 9281
rect 12137 9255 12138 9281
rect 12110 8834 12138 9255
rect 12334 9282 12362 9590
rect 12334 9249 12362 9254
rect 12726 10009 12754 10015
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12614 9226 12642 9231
rect 12614 9179 12642 9198
rect 12446 8946 12474 8951
rect 12446 8899 12474 8918
rect 12110 8801 12138 8806
rect 12446 8834 12474 8839
rect 12446 8787 12474 8806
rect 12726 8834 12754 9983
rect 12782 9954 12810 9959
rect 12782 9337 12810 9926
rect 12782 9311 12783 9337
rect 12809 9311 12810 9337
rect 12782 9305 12810 9311
rect 12726 8801 12754 8806
rect 12278 8778 12306 8783
rect 12278 8731 12306 8750
rect 11606 8409 11634 8414
rect 12670 8386 12698 8391
rect 11494 8073 11522 8078
rect 12334 8105 12362 8111
rect 12334 8079 12335 8105
rect 12361 8079 12362 8105
rect 10934 8050 10962 8055
rect 10262 8022 10458 8050
rect 10878 8049 10962 8050
rect 10878 8023 10935 8049
rect 10961 8023 10962 8049
rect 10878 8022 10962 8023
rect 10262 7993 10290 8022
rect 10262 7967 10263 7993
rect 10289 7967 10290 7993
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9254 7713 9282 7719
rect 9254 7687 9255 7713
rect 9281 7687 9282 7713
rect 9086 7658 9114 7663
rect 9086 7611 9114 7630
rect 9142 7657 9170 7663
rect 9142 7631 9143 7657
rect 9169 7631 9170 7657
rect 9030 6847 9031 6873
rect 9057 6847 9058 6873
rect 9030 6841 9058 6847
rect 9142 6762 9170 7631
rect 9198 7321 9226 7327
rect 9198 7295 9199 7321
rect 9225 7295 9226 7321
rect 9198 7154 9226 7295
rect 9198 7121 9226 7126
rect 8918 6734 9170 6762
rect 8134 6511 8135 6537
rect 8161 6511 8162 6537
rect 8134 6505 8162 6511
rect 9198 6538 9226 6543
rect 9254 6538 9282 7687
rect 9310 7657 9338 7663
rect 9310 7631 9311 7657
rect 9337 7631 9338 7657
rect 9310 7322 9338 7631
rect 9422 7658 9450 7663
rect 9422 7377 9450 7630
rect 9422 7351 9423 7377
rect 9449 7351 9450 7377
rect 9422 7345 9450 7351
rect 9310 7289 9338 7294
rect 9478 7322 9506 7327
rect 9198 6537 9282 6538
rect 9198 6511 9199 6537
rect 9225 6511 9282 6537
rect 9198 6510 9282 6511
rect 9366 7266 9394 7271
rect 9366 6538 9394 7238
rect 9478 7265 9506 7294
rect 9478 7239 9479 7265
rect 9505 7239 9506 7265
rect 9478 7233 9506 7239
rect 9702 7266 9730 7271
rect 9702 7219 9730 7238
rect 10150 7266 10178 7271
rect 10094 7209 10122 7215
rect 10094 7183 10095 7209
rect 10121 7183 10122 7209
rect 9422 7154 9450 7159
rect 9422 6986 9450 7126
rect 10094 7098 10122 7183
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10094 7065 10122 7070
rect 9918 7037 10050 7042
rect 10038 6986 10066 6991
rect 9422 6958 9674 6986
rect 9422 6538 9450 6543
rect 9366 6537 9450 6538
rect 9366 6511 9423 6537
rect 9449 6511 9450 6537
rect 9366 6510 9450 6511
rect 7798 6455 7799 6481
rect 7825 6455 7826 6481
rect 7798 6449 7826 6455
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 9030 1778 9058 1783
rect 9198 1778 9226 6510
rect 9422 6202 9450 6510
rect 9422 6201 9618 6202
rect 9422 6175 9423 6201
rect 9449 6175 9618 6201
rect 9422 6174 9618 6175
rect 9422 6169 9450 6174
rect 9590 6089 9618 6174
rect 9590 6063 9591 6089
rect 9617 6063 9618 6089
rect 9590 6057 9618 6063
rect 9646 2169 9674 6958
rect 9982 6958 10038 6986
rect 9982 6929 10010 6958
rect 10038 6953 10066 6958
rect 9982 6903 9983 6929
rect 10009 6903 10010 6929
rect 9982 6897 10010 6903
rect 10094 6929 10122 6935
rect 10094 6903 10095 6929
rect 10121 6903 10122 6929
rect 10094 6874 10122 6903
rect 10150 6929 10178 7238
rect 10262 7265 10290 7967
rect 10318 7938 10346 7943
rect 10318 7937 10402 7938
rect 10318 7911 10319 7937
rect 10345 7911 10402 7937
rect 10318 7910 10402 7911
rect 10318 7905 10346 7910
rect 10262 7239 10263 7265
rect 10289 7239 10290 7265
rect 10262 7233 10290 7239
rect 10318 7770 10346 7775
rect 10150 6903 10151 6929
rect 10177 6903 10178 6929
rect 10150 6897 10178 6903
rect 10206 7153 10234 7159
rect 10206 7127 10207 7153
rect 10233 7127 10234 7153
rect 10094 6841 10122 6846
rect 10206 6762 10234 7127
rect 10318 6873 10346 7742
rect 10374 7266 10402 7910
rect 10878 7770 10906 8022
rect 10934 8017 10962 8022
rect 11886 8050 11914 8055
rect 10878 7737 10906 7742
rect 11886 7769 11914 8022
rect 11886 7743 11887 7769
rect 11913 7743 11914 7769
rect 11886 7737 11914 7743
rect 12222 7938 12250 7943
rect 11998 7658 12026 7663
rect 11998 7657 12082 7658
rect 11998 7631 11999 7657
rect 12025 7631 12082 7657
rect 11998 7630 12082 7631
rect 11998 7625 12026 7630
rect 10990 7602 11018 7607
rect 10654 7266 10682 7271
rect 10374 7265 10682 7266
rect 10374 7239 10375 7265
rect 10401 7239 10655 7265
rect 10681 7239 10682 7265
rect 10374 7238 10682 7239
rect 10374 7233 10402 7238
rect 10654 7233 10682 7238
rect 10990 7265 11018 7574
rect 11830 7602 11858 7607
rect 11942 7601 11970 7607
rect 11942 7575 11943 7601
rect 11969 7575 11970 7601
rect 11942 7574 11970 7575
rect 11830 7546 11970 7574
rect 11998 7546 12026 7551
rect 10990 7239 10991 7265
rect 11017 7239 11018 7265
rect 10990 7233 11018 7239
rect 10766 7210 10794 7215
rect 10766 7163 10794 7182
rect 10822 7153 10850 7159
rect 10822 7127 10823 7153
rect 10849 7127 10850 7153
rect 10822 6986 10850 7127
rect 10710 6958 10850 6986
rect 11998 6986 12026 7518
rect 10710 6929 10738 6958
rect 11998 6939 12026 6958
rect 10710 6903 10711 6929
rect 10737 6903 10738 6929
rect 10710 6897 10738 6903
rect 10318 6847 10319 6873
rect 10345 6847 10346 6873
rect 10318 6841 10346 6847
rect 10094 6734 10234 6762
rect 11774 6818 11802 6823
rect 12054 6818 12082 7630
rect 12222 7657 12250 7910
rect 12334 7826 12362 8079
rect 12614 8106 12642 8111
rect 12502 8050 12530 8055
rect 12502 8003 12530 8022
rect 12558 8050 12586 8055
rect 12614 8050 12642 8078
rect 12558 8049 12642 8050
rect 12558 8023 12559 8049
rect 12585 8023 12642 8049
rect 12558 8022 12642 8023
rect 12558 8017 12586 8022
rect 12614 7937 12642 7943
rect 12614 7911 12615 7937
rect 12641 7911 12642 7937
rect 12614 7826 12642 7911
rect 12334 7798 12642 7826
rect 12222 7631 12223 7657
rect 12249 7631 12250 7657
rect 12222 7625 12250 7631
rect 12502 7714 12530 7719
rect 12502 7574 12530 7686
rect 12502 7546 12586 7574
rect 12558 7265 12586 7546
rect 12558 7239 12559 7265
rect 12585 7239 12586 7265
rect 12558 7233 12586 7239
rect 12614 7098 12642 7798
rect 12670 7826 12698 8358
rect 12782 8330 12810 8335
rect 12810 8302 12866 8330
rect 12782 8297 12810 8302
rect 12726 8050 12754 8055
rect 12754 8022 12810 8050
rect 12726 8017 12754 8022
rect 12726 7938 12754 7943
rect 12726 7891 12754 7910
rect 12670 7793 12698 7798
rect 12670 7714 12698 7719
rect 12782 7714 12810 8022
rect 12838 7769 12866 8302
rect 12838 7743 12839 7769
rect 12865 7743 12866 7769
rect 12838 7737 12866 7743
rect 12698 7686 12810 7714
rect 12670 7667 12698 7686
rect 12894 7574 12922 10262
rect 13230 10009 13258 10015
rect 13230 9983 13231 10009
rect 13257 9983 13258 10009
rect 13230 9954 13258 9983
rect 13230 9921 13258 9926
rect 13286 9953 13314 11159
rect 13342 10738 13370 11270
rect 13342 10705 13370 10710
rect 13286 9927 13287 9953
rect 13313 9927 13314 9953
rect 13286 9921 13314 9927
rect 13342 10346 13370 10351
rect 13342 10009 13370 10318
rect 13342 9983 13343 10009
rect 13369 9983 13370 10009
rect 13342 9338 13370 9983
rect 13398 9954 13426 11326
rect 13846 11186 13874 11191
rect 13790 10401 13818 10407
rect 13790 10375 13791 10401
rect 13817 10375 13818 10401
rect 13454 10066 13482 10071
rect 13454 10019 13482 10038
rect 13398 9921 13426 9926
rect 13622 10009 13650 10015
rect 13622 9983 13623 10009
rect 13649 9983 13650 10009
rect 13622 9730 13650 9983
rect 13734 10010 13762 10015
rect 13734 9963 13762 9982
rect 13454 9702 13650 9730
rect 13678 9953 13706 9959
rect 13678 9927 13679 9953
rect 13705 9927 13706 9953
rect 13454 9338 13482 9702
rect 13678 9674 13706 9927
rect 13286 9310 13370 9338
rect 13398 9310 13482 9338
rect 13510 9646 13706 9674
rect 12950 9282 12978 9287
rect 12950 8497 12978 9254
rect 13118 9282 13146 9287
rect 13286 9282 13314 9310
rect 13118 9281 13314 9282
rect 13118 9255 13119 9281
rect 13145 9255 13314 9281
rect 13118 9254 13314 9255
rect 13118 9249 13146 9254
rect 12950 8471 12951 8497
rect 12977 8471 12978 8497
rect 12950 8465 12978 8471
rect 13006 9225 13034 9231
rect 13006 9199 13007 9225
rect 13033 9199 13034 9225
rect 13006 8834 13034 9199
rect 13006 8049 13034 8806
rect 13006 8023 13007 8049
rect 13033 8023 13034 8049
rect 13006 8017 13034 8023
rect 13062 8441 13090 8447
rect 13062 8415 13063 8441
rect 13089 8415 13090 8441
rect 13062 8050 13090 8415
rect 13062 8017 13090 8022
rect 13118 7937 13146 7943
rect 13118 7911 13119 7937
rect 13145 7911 13146 7937
rect 13062 7770 13090 7775
rect 13062 7657 13090 7742
rect 13062 7631 13063 7657
rect 13089 7631 13090 7657
rect 13062 7625 13090 7631
rect 12782 7546 12922 7574
rect 12670 7266 12698 7271
rect 12782 7266 12810 7546
rect 12670 7265 12810 7266
rect 12670 7239 12671 7265
rect 12697 7239 12810 7265
rect 12670 7238 12810 7239
rect 13118 7266 13146 7911
rect 13174 7938 13202 9254
rect 13342 9225 13370 9231
rect 13342 9199 13343 9225
rect 13369 9199 13370 9225
rect 13342 8946 13370 9199
rect 13342 8913 13370 8918
rect 13230 8890 13258 8895
rect 13230 8834 13258 8862
rect 13398 8834 13426 9310
rect 13510 9281 13538 9646
rect 13510 9255 13511 9281
rect 13537 9255 13538 9281
rect 13510 9249 13538 9255
rect 13678 9561 13706 9567
rect 13678 9535 13679 9561
rect 13705 9535 13706 9561
rect 13678 9226 13706 9535
rect 13454 9170 13482 9175
rect 13454 9123 13482 9142
rect 13230 8806 13426 8834
rect 13230 8441 13258 8806
rect 13510 8721 13538 8727
rect 13510 8695 13511 8721
rect 13537 8695 13538 8721
rect 13230 8415 13231 8441
rect 13257 8415 13258 8441
rect 13230 8409 13258 8415
rect 13342 8553 13370 8559
rect 13342 8527 13343 8553
rect 13369 8527 13370 8553
rect 13230 8330 13258 8335
rect 13230 8283 13258 8302
rect 13174 7905 13202 7910
rect 13342 7714 13370 8527
rect 13510 8442 13538 8695
rect 13622 8442 13650 8447
rect 13678 8442 13706 9198
rect 13790 8834 13818 10375
rect 13846 10401 13874 11158
rect 14294 11073 14322 11079
rect 14294 11047 14295 11073
rect 14321 11047 14322 11073
rect 14294 10906 14322 11047
rect 14518 10906 14546 10911
rect 14322 10878 14378 10906
rect 14294 10873 14322 10878
rect 13958 10738 13986 10743
rect 13958 10457 13986 10710
rect 14294 10737 14322 10743
rect 14294 10711 14295 10737
rect 14321 10711 14322 10737
rect 14294 10682 14322 10711
rect 14294 10649 14322 10654
rect 14238 10514 14266 10519
rect 13958 10431 13959 10457
rect 13985 10431 13986 10457
rect 13958 10425 13986 10431
rect 14070 10513 14266 10514
rect 14070 10487 14239 10513
rect 14265 10487 14266 10513
rect 14070 10486 14266 10487
rect 13846 10375 13847 10401
rect 13873 10375 13874 10401
rect 13846 10369 13874 10375
rect 14070 10401 14098 10486
rect 14238 10481 14266 10486
rect 14070 10375 14071 10401
rect 14097 10375 14098 10401
rect 14070 10369 14098 10375
rect 14238 10402 14266 10407
rect 14182 10346 14210 10351
rect 14182 10299 14210 10318
rect 14238 10345 14266 10374
rect 14238 10319 14239 10345
rect 14265 10319 14266 10345
rect 14238 10313 14266 10319
rect 14350 10178 14378 10878
rect 14518 10794 14546 10878
rect 14798 10906 14826 12279
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 14798 10873 14826 10878
rect 18830 11185 18858 11191
rect 18830 11159 18831 11185
rect 18857 11159 18858 11185
rect 18830 10906 18858 11159
rect 18830 10873 18858 10878
rect 18830 10794 18858 10799
rect 14518 10793 14658 10794
rect 14518 10767 14519 10793
rect 14545 10767 14658 10793
rect 14518 10766 14658 10767
rect 14518 10761 14546 10766
rect 14238 10150 14378 10178
rect 14406 10682 14434 10687
rect 13846 10065 13874 10071
rect 13846 10039 13847 10065
rect 13873 10039 13874 10065
rect 13846 9954 13874 10039
rect 13846 9921 13874 9926
rect 14238 9226 14266 10150
rect 14406 10066 14434 10654
rect 14630 10457 14658 10766
rect 18830 10747 18858 10766
rect 20006 10794 20034 11215
rect 20006 10761 20034 10766
rect 14854 10738 14882 10743
rect 14854 10691 14882 10710
rect 15918 10737 15946 10743
rect 15918 10711 15919 10737
rect 15945 10711 15946 10737
rect 14630 10431 14631 10457
rect 14657 10431 14658 10457
rect 14630 10425 14658 10431
rect 15918 10682 15946 10711
rect 15918 10402 15946 10654
rect 20006 10681 20034 10687
rect 20006 10655 20007 10681
rect 20033 10655 20034 10681
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10458 20034 10655
rect 20006 10425 20034 10430
rect 15918 10369 15946 10374
rect 14406 10033 14434 10038
rect 14238 9193 14266 9198
rect 15134 10010 15162 10015
rect 15134 9618 15162 9982
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 14070 9170 14098 9175
rect 14070 9123 14098 9142
rect 15134 9169 15162 9590
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 15134 9143 15135 9169
rect 15161 9143 15162 9169
rect 15134 9137 15162 9143
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 14070 8946 14098 8951
rect 14070 8899 14098 8918
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 13958 8834 13986 8839
rect 13790 8833 13986 8834
rect 13790 8807 13959 8833
rect 13985 8807 13986 8833
rect 13790 8806 13986 8807
rect 13958 8610 13986 8806
rect 14182 8834 14210 8839
rect 14182 8787 14210 8806
rect 14630 8834 14658 8839
rect 14630 8787 14658 8806
rect 14742 8834 14770 8839
rect 14742 8787 14770 8806
rect 15246 8834 15274 8839
rect 14574 8777 14602 8783
rect 14574 8751 14575 8777
rect 14601 8751 14602 8777
rect 13958 8577 13986 8582
rect 14126 8721 14154 8727
rect 14126 8695 14127 8721
rect 14153 8695 14154 8721
rect 14126 8498 14154 8695
rect 14182 8498 14210 8503
rect 14126 8497 14210 8498
rect 14126 8471 14183 8497
rect 14209 8471 14210 8497
rect 14126 8470 14210 8471
rect 14182 8465 14210 8470
rect 13510 8414 13622 8442
rect 13650 8414 13706 8442
rect 13846 8442 13874 8461
rect 13622 8395 13650 8414
rect 13846 8409 13874 8414
rect 13790 8386 13818 8391
rect 13790 8161 13818 8358
rect 14574 8386 14602 8751
rect 14574 8353 14602 8358
rect 15246 8385 15274 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 15246 8359 15247 8385
rect 15273 8359 15274 8385
rect 15246 8353 15274 8359
rect 18830 8441 18858 8447
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 13790 8135 13791 8161
rect 13817 8135 13818 8161
rect 13790 8129 13818 8135
rect 13846 8330 13874 8335
rect 13846 8105 13874 8302
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 13846 8079 13847 8105
rect 13873 8079 13874 8105
rect 13846 8073 13874 8079
rect 13958 8049 13986 8055
rect 13958 8023 13959 8049
rect 13985 8023 13986 8049
rect 13454 7714 13482 7719
rect 13342 7713 13482 7714
rect 13342 7687 13455 7713
rect 13481 7687 13482 7713
rect 13342 7686 13482 7687
rect 13454 7681 13482 7686
rect 13958 7602 13986 8023
rect 13958 7569 13986 7574
rect 14294 7658 14322 7663
rect 12670 7233 12698 7238
rect 13118 7219 13146 7238
rect 12838 7210 12866 7215
rect 12950 7210 12978 7215
rect 12838 7209 12978 7210
rect 12838 7183 12839 7209
rect 12865 7183 12951 7209
rect 12977 7183 12978 7209
rect 12838 7182 12978 7183
rect 12838 7177 12866 7182
rect 12950 7177 12978 7182
rect 12782 7153 12810 7159
rect 12782 7127 12783 7153
rect 12809 7127 12810 7153
rect 12614 7070 12698 7098
rect 12614 6986 12642 6991
rect 12614 6873 12642 6958
rect 12614 6847 12615 6873
rect 12641 6847 12642 6873
rect 12614 6841 12642 6847
rect 11774 6817 12082 6818
rect 11774 6791 11775 6817
rect 11801 6791 12082 6817
rect 11774 6790 12082 6791
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 10094 6202 10122 6734
rect 9982 6174 10122 6202
rect 10878 6706 10906 6711
rect 9982 6145 10010 6174
rect 9982 6119 9983 6145
rect 10009 6119 10010 6145
rect 9982 6113 10010 6119
rect 10878 5922 10906 6678
rect 11046 6033 11074 6039
rect 11046 6007 11047 6033
rect 11073 6007 11074 6033
rect 11046 5922 11074 6007
rect 10878 5894 11074 5922
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9646 2143 9647 2169
rect 9673 2143 9674 2169
rect 9646 2137 9674 2143
rect 9422 2058 9450 2063
rect 9030 1777 9226 1778
rect 9030 1751 9031 1777
rect 9057 1751 9226 1777
rect 9030 1750 9226 1751
rect 9310 1833 9338 1839
rect 9310 1807 9311 1833
rect 9337 1807 9338 1833
rect 9030 1745 9058 1750
rect 9310 1694 9338 1807
rect 9086 1666 9338 1694
rect 9086 400 9114 1666
rect 9422 400 9450 2030
rect 10038 2058 10066 2063
rect 10038 2011 10066 2030
rect 10766 1834 10794 1839
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10766 400 10794 1806
rect 10878 1777 10906 5894
rect 11774 5362 11802 6790
rect 11774 5334 12194 5362
rect 12110 2058 12138 2063
rect 11214 1834 11242 1839
rect 11214 1787 11242 1806
rect 11774 1834 11802 1839
rect 10878 1751 10879 1777
rect 10905 1751 10906 1777
rect 10878 1745 10906 1751
rect 11774 400 11802 1806
rect 12110 400 12138 2030
rect 12166 1778 12194 5334
rect 12614 2170 12642 2175
rect 12670 2170 12698 7070
rect 12782 6986 12810 7127
rect 13062 7153 13090 7159
rect 13062 7127 13063 7153
rect 13089 7127 13090 7153
rect 12782 6958 13034 6986
rect 13006 6929 13034 6958
rect 13006 6903 13007 6929
rect 13033 6903 13034 6929
rect 13006 6897 13034 6903
rect 13062 6818 13090 7127
rect 14294 6985 14322 7630
rect 14742 7658 14770 7663
rect 14742 7611 14770 7630
rect 14518 7602 14546 7607
rect 14518 7555 14546 7574
rect 18830 7602 18858 8415
rect 20006 8329 20034 8335
rect 20006 8303 20007 8329
rect 20033 8303 20034 8329
rect 20006 8106 20034 8303
rect 20006 8073 20034 8078
rect 18830 7569 18858 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 14294 6959 14295 6985
rect 14321 6959 14322 6985
rect 14294 6953 14322 6959
rect 13062 6785 13090 6790
rect 14070 6818 14098 6823
rect 14070 4214 14098 6790
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 13958 4186 14098 4214
rect 12614 2169 12698 2170
rect 12614 2143 12615 2169
rect 12641 2143 12698 2169
rect 12614 2142 12698 2143
rect 13006 2617 13034 2623
rect 13006 2591 13007 2617
rect 13033 2591 13034 2617
rect 12614 2137 12642 2142
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1778 12306 1783
rect 12166 1777 12306 1778
rect 12166 1751 12279 1777
rect 12305 1751 12306 1777
rect 12166 1750 12306 1751
rect 12278 1745 12306 1750
rect 13006 1694 13034 2591
rect 13958 2561 13986 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 13958 2535 13959 2561
rect 13985 2535 13986 2561
rect 13958 2529 13986 2535
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12894 1666 13034 1694
rect 12894 490 12922 1666
rect 12782 462 12922 490
rect 12782 400 12810 462
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 10752 0 10808 400
rect 11760 0 11816 400
rect 12096 0 12152 400
rect 12768 0 12824 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8750 19110 8778 19138
rect 9310 19137 9338 19138
rect 9310 19111 9311 19137
rect 9311 19111 9337 19137
rect 9337 19111 9338 19137
rect 9310 19110 9338 19111
rect 8078 18718 8106 18746
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 8190 14182 8218 14210
rect 2086 13790 2114 13818
rect 966 12446 994 12474
rect 966 11465 994 11466
rect 966 11439 967 11465
rect 967 11439 993 11465
rect 993 11439 994 11465
rect 966 11438 994 11439
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 7350 13873 7378 13874
rect 7350 13847 7351 13873
rect 7351 13847 7377 13873
rect 7377 13847 7378 13873
rect 7350 13846 7378 13847
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2142 12753 2170 12754
rect 2142 12727 2143 12753
rect 2143 12727 2169 12753
rect 2169 12727 2170 12753
rect 2142 12726 2170 12727
rect 6510 12726 6538 12754
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9198 18745 9226 18746
rect 9198 18719 9199 18745
rect 9199 18719 9225 18745
rect 9225 18719 9226 18745
rect 9198 18718 9226 18719
rect 10766 19110 10794 19138
rect 11214 19137 11242 19138
rect 11214 19111 11215 19137
rect 11215 19111 11241 19137
rect 11241 19111 11242 19137
rect 11214 19110 11242 19111
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 11774 19110 11802 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 10094 18718 10122 18746
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 10710 18745 10738 18746
rect 10710 18719 10711 18745
rect 10711 18719 10737 18745
rect 10737 18719 10738 18745
rect 10710 18718 10738 18719
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 8694 14182 8722 14210
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9926 14265 9954 14266
rect 9926 14239 9927 14265
rect 9927 14239 9953 14265
rect 9953 14239 9954 14265
rect 9926 14238 9954 14239
rect 8806 14182 8834 14210
rect 8526 13846 8554 13874
rect 8022 13398 8050 13426
rect 7126 13342 7154 13370
rect 7574 13342 7602 13370
rect 7630 13118 7658 13146
rect 7014 12614 7042 12642
rect 6510 12222 6538 12250
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 8302 12809 8330 12810
rect 8302 12783 8303 12809
rect 8303 12783 8329 12809
rect 8329 12783 8330 12809
rect 8302 12782 8330 12783
rect 7966 12614 7994 12642
rect 8246 12614 8274 12642
rect 7742 11969 7770 11970
rect 7742 11943 7743 11969
rect 7743 11943 7769 11969
rect 7769 11943 7770 11969
rect 7742 11942 7770 11943
rect 8246 12222 8274 12250
rect 7966 11774 7994 11802
rect 2142 11577 2170 11578
rect 2142 11551 2143 11577
rect 2143 11551 2169 11577
rect 2169 11551 2170 11577
rect 2142 11550 2170 11551
rect 5894 11550 5922 11578
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 7350 11494 7378 11522
rect 7574 11633 7602 11634
rect 7574 11607 7575 11633
rect 7575 11607 7601 11633
rect 7601 11607 7602 11633
rect 7574 11606 7602 11607
rect 7574 11494 7602 11522
rect 7742 11577 7770 11578
rect 7742 11551 7743 11577
rect 7743 11551 7769 11577
rect 7769 11551 7770 11577
rect 7742 11550 7770 11551
rect 7910 11577 7938 11578
rect 7910 11551 7911 11577
rect 7911 11551 7937 11577
rect 7937 11551 7938 11577
rect 7910 11550 7938 11551
rect 8190 11942 8218 11970
rect 8526 13398 8554 13426
rect 9086 13873 9114 13874
rect 9086 13847 9087 13873
rect 9087 13847 9113 13873
rect 9113 13847 9114 13873
rect 9086 13846 9114 13847
rect 9478 13873 9506 13874
rect 9478 13847 9479 13873
rect 9479 13847 9505 13873
rect 9505 13847 9506 13873
rect 9478 13846 9506 13847
rect 8806 13398 8834 13426
rect 8694 13174 8722 13202
rect 8974 13201 9002 13202
rect 8974 13175 8975 13201
rect 8975 13175 9001 13201
rect 9001 13175 9002 13201
rect 8974 13174 9002 13175
rect 10318 14265 10346 14266
rect 10318 14239 10319 14265
rect 10319 14239 10345 14265
rect 10345 14239 10346 14265
rect 10318 14238 10346 14239
rect 11046 14238 11074 14266
rect 9982 14182 10010 14210
rect 10374 14182 10402 14210
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9814 13201 9842 13202
rect 9814 13175 9815 13201
rect 9815 13175 9841 13201
rect 9841 13175 9842 13201
rect 9814 13174 9842 13175
rect 10262 13201 10290 13202
rect 10262 13175 10263 13201
rect 10263 13175 10289 13201
rect 10289 13175 10290 13201
rect 10262 13174 10290 13175
rect 10654 13174 10682 13202
rect 9086 13145 9114 13146
rect 9086 13119 9087 13145
rect 9087 13119 9113 13145
rect 9113 13119 9114 13145
rect 9086 13118 9114 13119
rect 8750 12782 8778 12810
rect 8694 12641 8722 12642
rect 8694 12615 8695 12641
rect 8695 12615 8721 12641
rect 8721 12615 8722 12641
rect 8694 12614 8722 12615
rect 9366 12614 9394 12642
rect 8358 12334 8386 12362
rect 8694 12361 8722 12362
rect 8694 12335 8695 12361
rect 8695 12335 8721 12361
rect 8721 12335 8722 12361
rect 8694 12334 8722 12335
rect 8470 12110 8498 12138
rect 8806 12110 8834 12138
rect 8918 11774 8946 11802
rect 8078 11550 8106 11578
rect 8134 11438 8162 11466
rect 7462 11073 7490 11074
rect 7462 11047 7463 11073
rect 7463 11047 7489 11073
rect 7489 11047 7490 11073
rect 7462 11046 7490 11047
rect 7574 11102 7602 11130
rect 7182 10793 7210 10794
rect 7182 10767 7183 10793
rect 7183 10767 7209 10793
rect 7209 10767 7210 10793
rect 7182 10766 7210 10767
rect 7574 10766 7602 10794
rect 6230 10710 6258 10738
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2086 10374 2114 10402
rect 6846 10737 6874 10738
rect 6846 10711 6847 10737
rect 6847 10711 6873 10737
rect 6873 10711 6874 10737
rect 6846 10710 6874 10711
rect 7070 10430 7098 10458
rect 7238 10401 7266 10402
rect 7238 10375 7239 10401
rect 7239 10375 7265 10401
rect 7265 10375 7266 10401
rect 7238 10374 7266 10375
rect 6006 10150 6034 10178
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 5614 9225 5642 9226
rect 5614 9199 5615 9225
rect 5615 9199 5641 9225
rect 5641 9199 5642 9225
rect 5614 9198 5642 9199
rect 7070 10150 7098 10178
rect 7406 10094 7434 10122
rect 8246 11102 8274 11130
rect 7910 10710 7938 10738
rect 7854 10374 7882 10402
rect 7518 9953 7546 9954
rect 7518 9927 7519 9953
rect 7519 9927 7545 9953
rect 7545 9927 7546 9953
rect 7518 9926 7546 9927
rect 7518 9561 7546 9562
rect 7518 9535 7519 9561
rect 7519 9535 7545 9561
rect 7545 9535 7546 9561
rect 7518 9534 7546 9535
rect 6790 9198 6818 9226
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 6734 8414 6762 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 966 8078 994 8106
rect 7014 9198 7042 9226
rect 7070 9478 7098 9506
rect 7406 9505 7434 9506
rect 7406 9479 7407 9505
rect 7407 9479 7433 9505
rect 7433 9479 7434 9505
rect 7406 9478 7434 9479
rect 8190 10710 8218 10738
rect 8526 11606 8554 11634
rect 8414 10262 8442 10290
rect 8078 10065 8106 10066
rect 8078 10039 8079 10065
rect 8079 10039 8105 10065
rect 8105 10039 8106 10065
rect 8078 10038 8106 10039
rect 7966 9982 7994 10010
rect 8302 10009 8330 10010
rect 8302 9983 8303 10009
rect 8303 9983 8329 10009
rect 8329 9983 8330 10009
rect 8302 9982 8330 9983
rect 8022 9953 8050 9954
rect 8022 9927 8023 9953
rect 8023 9927 8049 9953
rect 8049 9927 8050 9953
rect 8022 9926 8050 9927
rect 7854 9870 7882 9898
rect 8358 9702 8386 9730
rect 7686 9478 7714 9506
rect 8358 9478 8386 9506
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 10990 12753 11018 12754
rect 10990 12727 10991 12753
rect 10991 12727 11017 12753
rect 11017 12727 11018 12753
rect 10990 12726 11018 12727
rect 11942 12726 11970 12754
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10542 12558 10570 12586
rect 10022 12530 10050 12531
rect 9814 12334 9842 12362
rect 9590 11942 9618 11970
rect 9478 11913 9506 11914
rect 9478 11887 9479 11913
rect 9479 11887 9505 11913
rect 9505 11887 9506 11913
rect 9478 11886 9506 11887
rect 9926 12110 9954 12138
rect 9814 11886 9842 11914
rect 9478 11774 9506 11802
rect 9702 11662 9730 11690
rect 8470 9422 8498 9450
rect 8414 9310 8442 9338
rect 8750 11438 8778 11466
rect 8638 10009 8666 10010
rect 8638 9983 8639 10009
rect 8639 9983 8665 10009
rect 8665 9983 8666 10009
rect 8638 9982 8666 9983
rect 7294 9225 7322 9226
rect 7294 9199 7295 9225
rect 7295 9199 7321 9225
rect 7321 9199 7322 9225
rect 7294 9198 7322 9199
rect 8526 9198 8554 9226
rect 8190 8806 8218 8834
rect 7126 8694 7154 8722
rect 7798 8526 7826 8554
rect 6734 8105 6762 8106
rect 6734 8079 6735 8105
rect 6735 8079 6761 8105
rect 6761 8079 6762 8105
rect 6734 8078 6762 8079
rect 8358 8721 8386 8722
rect 8358 8695 8359 8721
rect 8359 8695 8385 8721
rect 8385 8695 8386 8721
rect 8358 8694 8386 8695
rect 8582 9702 8610 9730
rect 8974 10038 9002 10066
rect 8862 9758 8890 9786
rect 8806 9310 8834 9338
rect 8750 9281 8778 9282
rect 8750 9255 8751 9281
rect 8751 9255 8777 9281
rect 8777 9255 8778 9281
rect 8750 9254 8778 9255
rect 8638 9142 8666 9170
rect 8694 9198 8722 9226
rect 8638 8862 8666 8890
rect 8470 8721 8498 8722
rect 8470 8695 8471 8721
rect 8471 8695 8497 8721
rect 8497 8695 8498 8721
rect 8470 8694 8498 8695
rect 8358 8049 8386 8050
rect 8358 8023 8359 8049
rect 8359 8023 8385 8049
rect 8385 8023 8386 8049
rect 8358 8022 8386 8023
rect 8134 7574 8162 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 7798 7265 7826 7266
rect 7798 7239 7799 7265
rect 7799 7239 7825 7265
rect 7825 7239 7826 7265
rect 7798 7238 7826 7239
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 8246 7238 8274 7266
rect 8526 8078 8554 8106
rect 8750 8833 8778 8834
rect 8750 8807 8751 8833
rect 8751 8807 8777 8833
rect 8777 8807 8778 8833
rect 8750 8806 8778 8807
rect 8862 8777 8890 8778
rect 8862 8751 8863 8777
rect 8863 8751 8889 8777
rect 8889 8751 8890 8777
rect 8862 8750 8890 8751
rect 8694 8553 8722 8554
rect 8694 8527 8695 8553
rect 8695 8527 8721 8553
rect 8721 8527 8722 8553
rect 8694 8526 8722 8527
rect 8806 8470 8834 8498
rect 9198 11633 9226 11634
rect 9198 11607 9199 11633
rect 9199 11607 9225 11633
rect 9225 11607 9226 11633
rect 9198 11606 9226 11607
rect 9758 11606 9786 11634
rect 9142 11158 9170 11186
rect 9366 11073 9394 11074
rect 9366 11047 9367 11073
rect 9367 11047 9393 11073
rect 9393 11047 9394 11073
rect 9366 11046 9394 11047
rect 9478 10542 9506 10570
rect 9702 11577 9730 11578
rect 9702 11551 9703 11577
rect 9703 11551 9729 11577
rect 9729 11551 9730 11577
rect 9702 11550 9730 11551
rect 9590 11185 9618 11186
rect 9590 11159 9591 11185
rect 9591 11159 9617 11185
rect 9617 11159 9618 11185
rect 9590 11158 9618 11159
rect 10150 12361 10178 12362
rect 10150 12335 10151 12361
rect 10151 12335 10177 12361
rect 10177 12335 10178 12361
rect 10150 12334 10178 12335
rect 10542 12110 10570 12138
rect 10038 11830 10066 11858
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9870 11662 9898 11690
rect 10262 11857 10290 11858
rect 10262 11831 10263 11857
rect 10263 11831 10289 11857
rect 10289 11831 10290 11857
rect 10262 11830 10290 11831
rect 10094 11633 10122 11634
rect 10094 11607 10095 11633
rect 10095 11607 10121 11633
rect 10121 11607 10122 11633
rect 10094 11606 10122 11607
rect 9926 11494 9954 11522
rect 10318 11438 10346 11466
rect 10318 11158 10346 11186
rect 10878 12641 10906 12642
rect 10878 12615 10879 12641
rect 10879 12615 10905 12641
rect 10905 12615 10906 12641
rect 10878 12614 10906 12615
rect 10766 11942 10794 11970
rect 11270 12558 11298 12586
rect 12222 12558 12250 12586
rect 12782 12558 12810 12586
rect 12782 12390 12810 12418
rect 12838 12222 12866 12250
rect 12446 12054 12474 12082
rect 12782 12054 12810 12082
rect 12670 12025 12698 12026
rect 12670 11999 12671 12025
rect 12671 11999 12697 12025
rect 12697 11999 12698 12025
rect 12670 11998 12698 11999
rect 11550 11942 11578 11970
rect 10934 11718 10962 11746
rect 10654 11550 10682 11578
rect 10374 11494 10402 11522
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9534 10766 9562 10794
rect 9198 9870 9226 9898
rect 9254 9534 9282 9562
rect 9478 9478 9506 9506
rect 9142 9422 9170 9450
rect 8974 9169 9002 9170
rect 8974 9143 8975 9169
rect 8975 9143 9001 9169
rect 9001 9143 9002 9169
rect 8974 9142 9002 9143
rect 9030 8918 9058 8946
rect 9086 9086 9114 9114
rect 8974 8721 9002 8722
rect 8974 8695 8975 8721
rect 8975 8695 9001 8721
rect 9001 8695 9002 8721
rect 8974 8694 9002 8695
rect 9254 9225 9282 9226
rect 9254 9199 9255 9225
rect 9255 9199 9281 9225
rect 9281 9199 9282 9225
rect 9254 9198 9282 9199
rect 9422 9198 9450 9226
rect 9590 9926 9618 9954
rect 9702 9702 9730 9730
rect 10094 10654 10122 10682
rect 10038 10318 10066 10346
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10206 10038 10234 10066
rect 10206 9729 10234 9730
rect 10206 9703 10207 9729
rect 10207 9703 10233 9729
rect 10233 9703 10234 9729
rect 10206 9702 10234 9703
rect 9534 9281 9562 9282
rect 9534 9255 9535 9281
rect 9535 9255 9561 9281
rect 9561 9255 9562 9281
rect 9534 9254 9562 9255
rect 9870 9561 9898 9562
rect 9870 9535 9871 9561
rect 9871 9535 9897 9561
rect 9897 9535 9898 9561
rect 9870 9534 9898 9535
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10262 9310 10290 9338
rect 10150 9254 10178 9282
rect 9814 9198 9842 9226
rect 10038 9225 10066 9226
rect 10038 9199 10039 9225
rect 10039 9199 10065 9225
rect 10065 9199 10066 9225
rect 10038 9198 10066 9199
rect 10262 8918 10290 8946
rect 9478 8833 9506 8834
rect 9478 8807 9479 8833
rect 9479 8807 9505 8833
rect 9505 8807 9506 8833
rect 9478 8806 9506 8807
rect 9086 8777 9114 8778
rect 9086 8751 9087 8777
rect 9087 8751 9113 8777
rect 9113 8751 9114 8777
rect 9086 8750 9114 8751
rect 10654 11185 10682 11186
rect 10654 11159 10655 11185
rect 10655 11159 10681 11185
rect 10681 11159 10682 11185
rect 10654 11158 10682 11159
rect 10822 11577 10850 11578
rect 10822 11551 10823 11577
rect 10823 11551 10849 11577
rect 10849 11551 10850 11577
rect 10822 11550 10850 11551
rect 10934 11158 10962 11186
rect 11326 11550 11354 11578
rect 11102 11129 11130 11130
rect 11102 11103 11103 11129
rect 11103 11103 11129 11129
rect 11129 11103 11130 11129
rect 11102 11102 11130 11103
rect 10486 10793 10514 10794
rect 10486 10767 10487 10793
rect 10487 10767 10513 10793
rect 10513 10767 10514 10793
rect 10486 10766 10514 10767
rect 10766 10710 10794 10738
rect 10430 10654 10458 10682
rect 10430 10542 10458 10570
rect 10374 9534 10402 9562
rect 10542 10038 10570 10066
rect 10934 10401 10962 10402
rect 10934 10375 10935 10401
rect 10935 10375 10961 10401
rect 10961 10375 10962 10401
rect 10934 10374 10962 10375
rect 10990 9590 11018 9618
rect 10542 9281 10570 9282
rect 10542 9255 10543 9281
rect 10543 9255 10569 9281
rect 10569 9255 10570 9281
rect 10542 9254 10570 9255
rect 10374 9142 10402 9170
rect 10318 8750 10346 8778
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9254 8497 9282 8498
rect 9254 8471 9255 8497
rect 9255 8471 9281 8497
rect 9281 8471 9282 8497
rect 9254 8470 9282 8471
rect 9030 8414 9058 8442
rect 9534 8441 9562 8442
rect 9534 8415 9535 8441
rect 9535 8415 9561 8441
rect 9561 8415 9562 8441
rect 9534 8414 9562 8415
rect 8974 8358 9002 8386
rect 9030 8302 9058 8330
rect 8974 7601 9002 7602
rect 8974 7575 8975 7601
rect 8975 7575 9001 7601
rect 9001 7575 9002 7601
rect 8974 7574 9002 7575
rect 8470 7182 8498 7210
rect 8974 7182 9002 7210
rect 8134 6790 8162 6818
rect 8862 6817 8890 6818
rect 8862 6791 8863 6817
rect 8863 6791 8889 6817
rect 8889 6791 8890 6817
rect 8862 6790 8890 6791
rect 9422 8329 9450 8330
rect 9422 8303 9423 8329
rect 9423 8303 9449 8329
rect 9449 8303 9450 8329
rect 9422 8302 9450 8303
rect 10766 9225 10794 9226
rect 10766 9199 10767 9225
rect 10767 9199 10793 9225
rect 10793 9199 10794 9225
rect 10766 9198 10794 9199
rect 10766 8806 10794 8834
rect 10990 9198 11018 9226
rect 10878 9142 10906 9170
rect 10934 9086 10962 9114
rect 11102 9337 11130 9338
rect 11102 9311 11103 9337
rect 11103 9311 11129 9337
rect 11129 9311 11130 9337
rect 11102 9310 11130 9311
rect 11550 11577 11578 11578
rect 11550 11551 11551 11577
rect 11551 11551 11577 11577
rect 11577 11551 11578 11577
rect 11550 11550 11578 11551
rect 13062 12782 13090 12810
rect 13510 12809 13538 12810
rect 13510 12783 13511 12809
rect 13511 12783 13537 12809
rect 13537 12783 13538 12809
rect 13510 12782 13538 12783
rect 13342 12670 13370 12698
rect 13006 12390 13034 12418
rect 12894 11857 12922 11858
rect 12894 11831 12895 11857
rect 12895 11831 12921 11857
rect 12921 11831 12922 11857
rect 12894 11830 12922 11831
rect 12782 11774 12810 11802
rect 13118 12222 13146 12250
rect 11886 11577 11914 11578
rect 11886 11551 11887 11577
rect 11887 11551 11913 11577
rect 11913 11551 11914 11577
rect 11886 11550 11914 11551
rect 12558 11577 12586 11578
rect 12558 11551 12559 11577
rect 12559 11551 12585 11577
rect 12585 11551 12586 11577
rect 12558 11550 12586 11551
rect 11886 11102 11914 11130
rect 11550 10374 11578 10402
rect 11382 10038 11410 10066
rect 10654 8582 10682 8610
rect 10934 8918 10962 8946
rect 11102 8833 11130 8834
rect 11102 8807 11103 8833
rect 11103 8807 11129 8833
rect 11129 8807 11130 8833
rect 11102 8806 11130 8807
rect 10654 8358 10682 8386
rect 10598 8302 10626 8330
rect 11494 8918 11522 8946
rect 11382 8889 11410 8890
rect 11382 8863 11383 8889
rect 11383 8863 11409 8889
rect 11409 8863 11410 8889
rect 11382 8862 11410 8863
rect 11382 8441 11410 8442
rect 11382 8415 11383 8441
rect 11383 8415 11409 8441
rect 11409 8415 11410 8441
rect 11382 8414 11410 8415
rect 11214 8358 11242 8386
rect 11158 8302 11186 8330
rect 11830 10822 11858 10850
rect 11662 9702 11690 9730
rect 11830 10345 11858 10346
rect 11830 10319 11831 10345
rect 11831 10319 11857 10345
rect 11857 10319 11858 10345
rect 11830 10318 11858 10319
rect 11774 10065 11802 10066
rect 11774 10039 11775 10065
rect 11775 10039 11801 10065
rect 11801 10039 11802 10065
rect 11774 10038 11802 10039
rect 11998 10849 12026 10850
rect 11998 10823 11999 10849
rect 11999 10823 12025 10849
rect 12025 10823 12026 10849
rect 11998 10822 12026 10823
rect 12278 10065 12306 10066
rect 12278 10039 12279 10065
rect 12279 10039 12305 10065
rect 12305 10039 12306 10065
rect 12278 10038 12306 10039
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 13790 12697 13818 12698
rect 13790 12671 13791 12697
rect 13791 12671 13817 12697
rect 13817 12671 13818 12697
rect 13790 12670 13818 12671
rect 13678 12558 13706 12586
rect 13398 12278 13426 12306
rect 14294 12697 14322 12698
rect 14294 12671 14295 12697
rect 14295 12671 14321 12697
rect 14321 12671 14322 12697
rect 14294 12670 14322 12671
rect 14182 12614 14210 12642
rect 14574 12641 14602 12642
rect 14574 12615 14575 12641
rect 14575 12615 14601 12641
rect 14601 12615 14602 12641
rect 14574 12614 14602 12615
rect 14742 12641 14770 12642
rect 14742 12615 14743 12641
rect 14743 12615 14769 12641
rect 14769 12615 14770 12641
rect 14742 12614 14770 12615
rect 18830 12753 18858 12754
rect 18830 12727 18831 12753
rect 18831 12727 18857 12753
rect 18857 12727 18858 12753
rect 18830 12726 18858 12727
rect 20006 13118 20034 13146
rect 19950 12782 19978 12810
rect 18942 12670 18970 12698
rect 18774 12614 18802 12642
rect 20006 12446 20034 12474
rect 18830 12361 18858 12362
rect 18830 12335 18831 12361
rect 18831 12335 18857 12361
rect 18857 12335 18858 12361
rect 18830 12334 18858 12335
rect 14518 12305 14546 12306
rect 14518 12279 14519 12305
rect 14519 12279 14545 12305
rect 14545 12279 14546 12305
rect 14518 12278 14546 12279
rect 13734 12110 13762 12138
rect 13286 11774 13314 11802
rect 13118 11185 13146 11186
rect 13118 11159 13119 11185
rect 13119 11159 13145 11185
rect 13145 11159 13146 11185
rect 13118 11158 13146 11159
rect 12838 10878 12866 10906
rect 12614 10065 12642 10066
rect 12614 10039 12615 10065
rect 12615 10039 12641 10065
rect 12641 10039 12642 10065
rect 12614 10038 12642 10039
rect 12894 10262 12922 10290
rect 12334 9590 12362 9618
rect 11942 9142 11970 9170
rect 12334 9254 12362 9282
rect 12614 9225 12642 9226
rect 12614 9199 12615 9225
rect 12615 9199 12641 9225
rect 12641 9199 12642 9225
rect 12614 9198 12642 9199
rect 12446 8945 12474 8946
rect 12446 8919 12447 8945
rect 12447 8919 12473 8945
rect 12473 8919 12474 8945
rect 12446 8918 12474 8919
rect 12110 8806 12138 8834
rect 12446 8833 12474 8834
rect 12446 8807 12447 8833
rect 12447 8807 12473 8833
rect 12473 8807 12474 8833
rect 12446 8806 12474 8807
rect 12782 9926 12810 9954
rect 12726 8806 12754 8834
rect 12278 8777 12306 8778
rect 12278 8751 12279 8777
rect 12279 8751 12305 8777
rect 12305 8751 12306 8777
rect 12278 8750 12306 8751
rect 11606 8414 11634 8442
rect 12670 8385 12698 8386
rect 12670 8359 12671 8385
rect 12671 8359 12697 8385
rect 12697 8359 12698 8385
rect 12670 8358 12698 8359
rect 11494 8078 11522 8106
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9086 7657 9114 7658
rect 9086 7631 9087 7657
rect 9087 7631 9113 7657
rect 9113 7631 9114 7657
rect 9086 7630 9114 7631
rect 9198 7126 9226 7154
rect 9422 7630 9450 7658
rect 9310 7294 9338 7322
rect 9478 7294 9506 7322
rect 9366 7238 9394 7266
rect 9702 7265 9730 7266
rect 9702 7239 9703 7265
rect 9703 7239 9729 7265
rect 9729 7239 9730 7265
rect 9702 7238 9730 7239
rect 10150 7238 10178 7266
rect 9422 7153 9450 7154
rect 9422 7127 9423 7153
rect 9423 7127 9449 7153
rect 9449 7127 9450 7153
rect 9422 7126 9450 7127
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10094 7070 10122 7098
rect 10022 7042 10050 7043
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 10038 6958 10066 6986
rect 10318 7742 10346 7770
rect 10094 6846 10122 6874
rect 11886 8022 11914 8050
rect 10878 7742 10906 7770
rect 12222 7910 12250 7938
rect 10990 7574 11018 7602
rect 11830 7574 11858 7602
rect 11998 7518 12026 7546
rect 10766 7209 10794 7210
rect 10766 7183 10767 7209
rect 10767 7183 10793 7209
rect 10793 7183 10794 7209
rect 10766 7182 10794 7183
rect 11998 6985 12026 6986
rect 11998 6959 11999 6985
rect 11999 6959 12025 6985
rect 12025 6959 12026 6985
rect 11998 6958 12026 6959
rect 12614 8078 12642 8106
rect 12502 8049 12530 8050
rect 12502 8023 12503 8049
rect 12503 8023 12529 8049
rect 12529 8023 12530 8049
rect 12502 8022 12530 8023
rect 12502 7686 12530 7714
rect 12782 8302 12810 8330
rect 12726 8022 12754 8050
rect 12726 7937 12754 7938
rect 12726 7911 12727 7937
rect 12727 7911 12753 7937
rect 12753 7911 12754 7937
rect 12726 7910 12754 7911
rect 12670 7798 12698 7826
rect 12670 7713 12698 7714
rect 12670 7687 12671 7713
rect 12671 7687 12697 7713
rect 12697 7687 12698 7713
rect 12670 7686 12698 7687
rect 13230 9926 13258 9954
rect 13342 10710 13370 10738
rect 13342 10318 13370 10346
rect 13846 11158 13874 11186
rect 13454 10065 13482 10066
rect 13454 10039 13455 10065
rect 13455 10039 13481 10065
rect 13481 10039 13482 10065
rect 13454 10038 13482 10039
rect 13398 9926 13426 9954
rect 13734 10009 13762 10010
rect 13734 9983 13735 10009
rect 13735 9983 13761 10009
rect 13761 9983 13762 10009
rect 13734 9982 13762 9983
rect 12950 9254 12978 9282
rect 13006 8806 13034 8834
rect 13062 8022 13090 8050
rect 13062 7742 13090 7770
rect 13342 8918 13370 8946
rect 13230 8862 13258 8890
rect 13678 9225 13706 9226
rect 13678 9199 13679 9225
rect 13679 9199 13705 9225
rect 13705 9199 13706 9225
rect 13678 9198 13706 9199
rect 13454 9169 13482 9170
rect 13454 9143 13455 9169
rect 13455 9143 13481 9169
rect 13481 9143 13482 9169
rect 13454 9142 13482 9143
rect 13230 8329 13258 8330
rect 13230 8303 13231 8329
rect 13231 8303 13257 8329
rect 13257 8303 13258 8329
rect 13230 8302 13258 8303
rect 13174 7910 13202 7938
rect 14294 10878 14322 10906
rect 13958 10710 13986 10738
rect 14294 10654 14322 10682
rect 14238 10374 14266 10402
rect 14182 10345 14210 10346
rect 14182 10319 14183 10345
rect 14183 10319 14209 10345
rect 14209 10319 14210 10345
rect 14182 10318 14210 10319
rect 14518 10878 14546 10906
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20006 12110 20034 12138
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 20006 11774 20034 11802
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14798 10878 14826 10906
rect 18830 10878 18858 10906
rect 14406 10654 14434 10682
rect 13846 9926 13874 9954
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20006 10766 20034 10794
rect 14854 10737 14882 10738
rect 14854 10711 14855 10737
rect 14855 10711 14881 10737
rect 14881 10711 14882 10737
rect 14854 10710 14882 10711
rect 15918 10654 15946 10682
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 20006 10430 20034 10458
rect 15918 10374 15946 10402
rect 14406 10038 14434 10066
rect 14238 9198 14266 9226
rect 15134 9982 15162 10010
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 15134 9590 15162 9618
rect 14070 9169 14098 9170
rect 14070 9143 14071 9169
rect 14071 9143 14097 9169
rect 14097 9143 14098 9169
rect 14070 9142 14098 9143
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 20006 9422 20034 9450
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14070 8945 14098 8946
rect 14070 8919 14071 8945
rect 14071 8919 14097 8945
rect 14097 8919 14098 8945
rect 14070 8918 14098 8919
rect 14182 8833 14210 8834
rect 14182 8807 14183 8833
rect 14183 8807 14209 8833
rect 14209 8807 14210 8833
rect 14182 8806 14210 8807
rect 14630 8833 14658 8834
rect 14630 8807 14631 8833
rect 14631 8807 14657 8833
rect 14657 8807 14658 8833
rect 14630 8806 14658 8807
rect 14742 8833 14770 8834
rect 14742 8807 14743 8833
rect 14743 8807 14769 8833
rect 14769 8807 14770 8833
rect 14742 8806 14770 8807
rect 15246 8806 15274 8834
rect 13958 8582 13986 8610
rect 13622 8441 13650 8442
rect 13622 8415 13623 8441
rect 13623 8415 13649 8441
rect 13649 8415 13650 8441
rect 13622 8414 13650 8415
rect 13846 8441 13874 8442
rect 13846 8415 13847 8441
rect 13847 8415 13873 8441
rect 13873 8415 13874 8441
rect 13846 8414 13874 8415
rect 13790 8358 13818 8386
rect 14574 8358 14602 8386
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 13846 8302 13874 8330
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 13958 7574 13986 7602
rect 14294 7630 14322 7658
rect 13118 7265 13146 7266
rect 13118 7239 13119 7265
rect 13119 7239 13145 7265
rect 13145 7239 13146 7265
rect 13118 7238 13146 7239
rect 12614 6958 12642 6986
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 10878 6678 10906 6706
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9422 2030 9450 2058
rect 10038 2057 10066 2058
rect 10038 2031 10039 2057
rect 10039 2031 10065 2057
rect 10065 2031 10066 2057
rect 10038 2030 10066 2031
rect 10766 1806 10794 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 12110 2030 12138 2058
rect 11214 1833 11242 1834
rect 11214 1807 11215 1833
rect 11215 1807 11241 1833
rect 11241 1807 11242 1833
rect 11214 1806 11242 1807
rect 11774 1806 11802 1834
rect 14742 7657 14770 7658
rect 14742 7631 14743 7657
rect 14743 7631 14769 7657
rect 14769 7631 14770 7657
rect 14742 7630 14770 7631
rect 14518 7601 14546 7602
rect 14518 7575 14519 7601
rect 14519 7575 14545 7601
rect 14545 7575 14546 7601
rect 14518 7574 14546 7575
rect 20006 8078 20034 8106
rect 18830 7574 18858 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 13062 6790 13090 6818
rect 14070 6817 14098 6818
rect 14070 6791 14071 6817
rect 14071 6791 14097 6817
rect 14097 6791 14098 6817
rect 14070 6790 14098 6791
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8745 19110 8750 19138
rect 8778 19110 9310 19138
rect 9338 19110 9343 19138
rect 10761 19110 10766 19138
rect 10794 19110 11214 19138
rect 11242 19110 11247 19138
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8073 18718 8078 18746
rect 8106 18718 9198 18746
rect 9226 18718 9231 18746
rect 10089 18718 10094 18746
rect 10122 18718 10710 18746
rect 10738 18718 10743 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9921 14238 9926 14266
rect 9954 14238 10094 14266
rect 10313 14238 10318 14266
rect 10346 14238 11046 14266
rect 11074 14238 11079 14266
rect 10066 14210 10094 14238
rect 8185 14182 8190 14210
rect 8218 14182 8694 14210
rect 8722 14182 8727 14210
rect 8801 14182 8806 14210
rect 8834 14182 9982 14210
rect 10010 14182 10015 14210
rect 10066 14182 10374 14210
rect 10402 14182 10407 14210
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 7345 13846 7350 13874
rect 7378 13846 8526 13874
rect 8554 13846 8559 13874
rect 9081 13846 9086 13874
rect 9114 13846 9478 13874
rect 9506 13846 9511 13874
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 8017 13398 8022 13426
rect 8050 13398 8526 13426
rect 8554 13398 8806 13426
rect 8834 13398 8839 13426
rect 7121 13342 7126 13370
rect 7154 13342 7574 13370
rect 7602 13342 7607 13370
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 8689 13174 8694 13202
rect 8722 13174 8974 13202
rect 9002 13174 9814 13202
rect 9842 13174 10262 13202
rect 10290 13174 10654 13202
rect 10682 13174 10687 13202
rect 20600 13146 21000 13160
rect 7625 13118 7630 13146
rect 7658 13118 9086 13146
rect 9114 13118 9119 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 20600 12810 21000 12824
rect 8297 12782 8302 12810
rect 8330 12782 8750 12810
rect 8778 12782 8783 12810
rect 13057 12782 13062 12810
rect 13090 12782 13510 12810
rect 13538 12782 15974 12810
rect 19945 12782 19950 12810
rect 19978 12782 21000 12810
rect 15946 12754 15974 12782
rect 20600 12768 21000 12782
rect 2137 12726 2142 12754
rect 2170 12726 6510 12754
rect 6538 12726 6543 12754
rect 10985 12726 10990 12754
rect 11018 12726 11942 12754
rect 11970 12726 11975 12754
rect 15946 12726 18830 12754
rect 18858 12726 18863 12754
rect 13337 12670 13342 12698
rect 13370 12670 13790 12698
rect 13818 12670 13823 12698
rect 14289 12670 14294 12698
rect 14322 12670 18942 12698
rect 18970 12670 18975 12698
rect 7009 12614 7014 12642
rect 7042 12614 7966 12642
rect 7994 12614 7999 12642
rect 8241 12614 8246 12642
rect 8274 12614 8694 12642
rect 8722 12614 9366 12642
rect 9394 12614 10878 12642
rect 10906 12614 10911 12642
rect 14177 12614 14182 12642
rect 14210 12614 14574 12642
rect 14602 12614 14607 12642
rect 14737 12614 14742 12642
rect 14770 12614 18774 12642
rect 18802 12614 18807 12642
rect 10537 12558 10542 12586
rect 10570 12558 11270 12586
rect 11298 12558 12222 12586
rect 12250 12558 12782 12586
rect 12810 12558 13678 12586
rect 13706 12558 13711 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 0 12474 400 12488
rect 20600 12474 21000 12488
rect 0 12446 966 12474
rect 994 12446 999 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 0 12432 400 12446
rect 20600 12432 21000 12446
rect 12777 12390 12782 12418
rect 12810 12390 13006 12418
rect 13034 12390 13039 12418
rect 8353 12334 8358 12362
rect 8386 12334 8694 12362
rect 8722 12334 9814 12362
rect 9842 12334 10150 12362
rect 10178 12334 10183 12362
rect 15946 12334 18830 12362
rect 18858 12334 18863 12362
rect 15946 12306 15974 12334
rect 13393 12278 13398 12306
rect 13426 12278 14518 12306
rect 14546 12278 15974 12306
rect 6505 12222 6510 12250
rect 6538 12222 8246 12250
rect 8274 12222 8279 12250
rect 12833 12222 12838 12250
rect 12866 12222 13118 12250
rect 13146 12222 13151 12250
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 8465 12110 8470 12138
rect 8498 12110 8806 12138
rect 8834 12110 9926 12138
rect 9954 12110 10542 12138
rect 10570 12110 13734 12138
rect 13762 12110 13767 12138
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 12441 12054 12446 12082
rect 12474 12054 12782 12082
rect 12810 12054 12815 12082
rect 12665 11998 12670 12026
rect 12698 11998 15974 12026
rect 15946 11970 15974 11998
rect 7737 11942 7742 11970
rect 7770 11942 8190 11970
rect 8218 11942 8223 11970
rect 9585 11942 9590 11970
rect 9618 11942 10766 11970
rect 10794 11942 11550 11970
rect 11578 11942 11583 11970
rect 15946 11942 18830 11970
rect 18858 11942 18863 11970
rect 9473 11886 9478 11914
rect 9506 11886 9814 11914
rect 9842 11886 9847 11914
rect 10033 11830 10038 11858
rect 10066 11830 10122 11858
rect 10257 11830 10262 11858
rect 10290 11830 12894 11858
rect 12922 11830 12927 11858
rect 7961 11774 7966 11802
rect 7994 11774 7999 11802
rect 8913 11774 8918 11802
rect 8946 11774 9478 11802
rect 9506 11774 9511 11802
rect 7966 11634 7994 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 10094 11746 10122 11830
rect 20600 11802 21000 11816
rect 12777 11774 12782 11802
rect 12810 11774 13286 11802
rect 13314 11774 13319 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 20600 11760 21000 11774
rect 10094 11718 10934 11746
rect 10962 11718 10967 11746
rect 9697 11662 9702 11690
rect 9730 11662 9870 11690
rect 9898 11662 9903 11690
rect 7569 11606 7574 11634
rect 7602 11606 8526 11634
rect 8554 11606 8559 11634
rect 9193 11606 9198 11634
rect 9226 11606 9758 11634
rect 9786 11606 10094 11634
rect 10122 11606 10127 11634
rect 2137 11550 2142 11578
rect 2170 11550 5894 11578
rect 5922 11550 7742 11578
rect 7770 11550 7775 11578
rect 7905 11550 7910 11578
rect 7938 11550 8078 11578
rect 8106 11550 8111 11578
rect 9697 11550 9702 11578
rect 9730 11550 10654 11578
rect 10682 11550 10687 11578
rect 10817 11550 10822 11578
rect 10850 11550 11326 11578
rect 11354 11550 11550 11578
rect 11578 11550 11583 11578
rect 11881 11550 11886 11578
rect 11914 11550 12558 11578
rect 12586 11550 12591 11578
rect 7345 11494 7350 11522
rect 7378 11494 7574 11522
rect 7602 11494 7607 11522
rect 9921 11494 9926 11522
rect 9954 11494 10374 11522
rect 10402 11494 10407 11522
rect 0 11466 400 11480
rect 0 11438 966 11466
rect 994 11438 999 11466
rect 8129 11438 8134 11466
rect 8162 11438 8750 11466
rect 8778 11438 10318 11466
rect 10346 11438 10351 11466
rect 0 11424 400 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9137 11158 9142 11186
rect 9170 11158 9590 11186
rect 9618 11158 9623 11186
rect 10313 11158 10318 11186
rect 10346 11158 10654 11186
rect 10682 11158 10687 11186
rect 10929 11158 10934 11186
rect 10962 11158 13118 11186
rect 13146 11158 13846 11186
rect 13874 11158 13879 11186
rect 7569 11102 7574 11130
rect 7602 11102 8246 11130
rect 8274 11102 11102 11130
rect 11130 11102 11886 11130
rect 11914 11102 11919 11130
rect 7457 11046 7462 11074
rect 7490 11046 9366 11074
rect 9394 11046 9399 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 12833 10878 12838 10906
rect 12866 10878 14294 10906
rect 14322 10878 14518 10906
rect 14546 10878 14798 10906
rect 14826 10878 14831 10906
rect 15946 10878 18830 10906
rect 18858 10878 18863 10906
rect 11825 10822 11830 10850
rect 11858 10822 11998 10850
rect 12026 10822 12031 10850
rect 7177 10766 7182 10794
rect 7210 10766 7574 10794
rect 7602 10766 7607 10794
rect 9529 10766 9534 10794
rect 9562 10766 10486 10794
rect 10514 10766 10519 10794
rect 15946 10738 15974 10878
rect 20600 10794 21000 10808
rect 18825 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 6225 10710 6230 10738
rect 6258 10710 6846 10738
rect 6874 10710 6879 10738
rect 7905 10710 7910 10738
rect 7938 10710 8190 10738
rect 8218 10710 10766 10738
rect 10794 10710 13342 10738
rect 13370 10710 13375 10738
rect 13953 10710 13958 10738
rect 13986 10710 14854 10738
rect 14882 10710 14887 10738
rect 14966 10710 15974 10738
rect 14966 10682 14994 10710
rect 18830 10682 18858 10766
rect 20600 10752 21000 10766
rect 10089 10654 10094 10682
rect 10122 10654 10430 10682
rect 10458 10654 10463 10682
rect 14289 10654 14294 10682
rect 14322 10654 14406 10682
rect 14434 10654 14994 10682
rect 15913 10654 15918 10682
rect 15946 10654 18858 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7546 10542 9478 10570
rect 9506 10542 10430 10570
rect 10458 10542 10463 10570
rect 7546 10458 7574 10542
rect 20600 10458 21000 10472
rect 7065 10430 7070 10458
rect 7098 10430 7574 10458
rect 20001 10430 20006 10458
rect 20034 10430 21000 10458
rect 20600 10416 21000 10430
rect 2081 10374 2086 10402
rect 2114 10374 4214 10402
rect 7233 10374 7238 10402
rect 7266 10374 7854 10402
rect 7882 10374 7887 10402
rect 9926 10374 10934 10402
rect 10962 10374 11550 10402
rect 11578 10374 11583 10402
rect 14233 10374 14238 10402
rect 14266 10374 15918 10402
rect 15946 10374 15951 10402
rect 4186 10346 4214 10374
rect 9926 10346 9954 10374
rect 4186 10318 9954 10346
rect 10033 10318 10038 10346
rect 10066 10318 11830 10346
rect 11858 10318 11863 10346
rect 13337 10318 13342 10346
rect 13370 10318 14182 10346
rect 14210 10318 14215 10346
rect 8409 10262 8414 10290
rect 8442 10262 12894 10290
rect 12922 10262 12927 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 6001 10150 6006 10178
rect 6034 10150 7070 10178
rect 7098 10150 7103 10178
rect 7401 10094 7406 10122
rect 7434 10094 10234 10122
rect 10206 10066 10234 10094
rect 8073 10038 8078 10066
rect 8106 10038 8974 10066
rect 9002 10038 9007 10066
rect 10201 10038 10206 10066
rect 10234 10038 10239 10066
rect 10537 10038 10542 10066
rect 10570 10038 11382 10066
rect 11410 10038 11774 10066
rect 11802 10038 11807 10066
rect 12273 10038 12278 10066
rect 12306 10038 12614 10066
rect 12642 10038 12647 10066
rect 13449 10038 13454 10066
rect 13482 10038 14406 10066
rect 14434 10038 14439 10066
rect 7961 9982 7966 10010
rect 7994 9982 8302 10010
rect 8330 9982 8638 10010
rect 8666 9982 8671 10010
rect 13729 9982 13734 10010
rect 13762 9982 15134 10010
rect 15162 9982 15167 10010
rect 7513 9926 7518 9954
rect 7546 9926 8022 9954
rect 8050 9926 9590 9954
rect 9618 9926 9623 9954
rect 12777 9926 12782 9954
rect 12810 9926 13230 9954
rect 13258 9926 13398 9954
rect 13426 9926 13846 9954
rect 13874 9926 13879 9954
rect 7849 9870 7854 9898
rect 7882 9870 9198 9898
rect 9226 9870 9231 9898
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 8843 9758 8862 9786
rect 8890 9758 8895 9786
rect 8353 9702 8358 9730
rect 8386 9702 8582 9730
rect 8610 9702 9702 9730
rect 9730 9702 9735 9730
rect 10201 9702 10206 9730
rect 10234 9702 11662 9730
rect 11690 9702 11695 9730
rect 10985 9590 10990 9618
rect 11018 9590 12334 9618
rect 12362 9590 12367 9618
rect 15129 9590 15134 9618
rect 15162 9590 18830 9618
rect 18858 9590 18863 9618
rect 7513 9534 7518 9562
rect 7546 9534 8386 9562
rect 9249 9534 9254 9562
rect 9282 9534 9870 9562
rect 9898 9534 10374 9562
rect 10402 9534 10407 9562
rect 8358 9506 8386 9534
rect 10990 9506 11018 9590
rect 7065 9478 7070 9506
rect 7098 9478 7406 9506
rect 7434 9478 7686 9506
rect 7714 9478 7719 9506
rect 8353 9478 8358 9506
rect 8386 9478 9478 9506
rect 9506 9478 9511 9506
rect 9590 9478 11018 9506
rect 9590 9450 9618 9478
rect 20600 9450 21000 9464
rect 8465 9422 8470 9450
rect 8498 9422 9142 9450
rect 9170 9422 9618 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 8395 9310 8414 9338
rect 8442 9310 8447 9338
rect 8801 9310 8806 9338
rect 8834 9310 10262 9338
rect 10290 9310 11102 9338
rect 11130 9310 11135 9338
rect 8745 9254 8750 9282
rect 8778 9254 9534 9282
rect 9562 9254 9567 9282
rect 10145 9254 10150 9282
rect 10178 9254 10542 9282
rect 10570 9254 10575 9282
rect 12329 9254 12334 9282
rect 12362 9254 12950 9282
rect 12978 9254 12983 9282
rect 5609 9198 5614 9226
rect 5642 9198 6790 9226
rect 6818 9198 7014 9226
rect 7042 9198 7294 9226
rect 7322 9198 8526 9226
rect 8554 9198 8559 9226
rect 8689 9198 8694 9226
rect 8722 9198 8862 9226
rect 8890 9198 8895 9226
rect 9249 9198 9254 9226
rect 9282 9198 9422 9226
rect 9450 9198 9814 9226
rect 9842 9198 9847 9226
rect 10033 9198 10038 9226
rect 10066 9198 10766 9226
rect 10794 9198 10799 9226
rect 10985 9198 10990 9226
rect 11018 9198 12614 9226
rect 12642 9198 12647 9226
rect 13673 9198 13678 9226
rect 13706 9198 14238 9226
rect 14266 9198 14271 9226
rect 8633 9142 8638 9170
rect 8666 9142 8974 9170
rect 9002 9142 9007 9170
rect 10369 9142 10374 9170
rect 10402 9142 10878 9170
rect 10906 9142 11942 9170
rect 11970 9142 11975 9170
rect 13449 9142 13454 9170
rect 13482 9142 14070 9170
rect 14098 9142 14103 9170
rect 9081 9086 9086 9114
rect 9114 9086 10934 9114
rect 10962 9086 10967 9114
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9025 8918 9030 8946
rect 9058 8918 10262 8946
rect 10290 8918 10934 8946
rect 10962 8918 11494 8946
rect 11522 8918 11527 8946
rect 12441 8918 12446 8946
rect 12474 8918 13342 8946
rect 13370 8918 14070 8946
rect 14098 8918 14103 8946
rect 8633 8862 8638 8890
rect 8666 8862 11382 8890
rect 11410 8862 13230 8890
rect 13258 8862 13263 8890
rect 8185 8806 8190 8834
rect 8218 8806 8750 8834
rect 8778 8806 9478 8834
rect 9506 8806 9511 8834
rect 10761 8806 10766 8834
rect 10794 8806 11102 8834
rect 11130 8806 11135 8834
rect 12105 8806 12110 8834
rect 12138 8806 12446 8834
rect 12474 8806 12726 8834
rect 12754 8806 13006 8834
rect 13034 8806 13039 8834
rect 14177 8806 14182 8834
rect 14210 8806 14630 8834
rect 14658 8806 14663 8834
rect 14737 8806 14742 8834
rect 14770 8806 15246 8834
rect 15274 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 8857 8750 8862 8778
rect 8890 8750 9086 8778
rect 9114 8750 9119 8778
rect 10313 8750 10318 8778
rect 10346 8750 12278 8778
rect 12306 8750 12311 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 7121 8694 7126 8722
rect 7154 8694 8358 8722
rect 8386 8694 8391 8722
rect 8465 8694 8470 8722
rect 8498 8694 8974 8722
rect 9002 8694 9007 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 10649 8582 10654 8610
rect 10682 8582 13958 8610
rect 13986 8582 13991 8610
rect 7793 8526 7798 8554
rect 7826 8526 8694 8554
rect 8722 8526 8727 8554
rect 8801 8470 8806 8498
rect 8834 8470 9254 8498
rect 9282 8470 9287 8498
rect 2137 8414 2142 8442
rect 2170 8414 6734 8442
rect 6762 8414 6767 8442
rect 9025 8414 9030 8442
rect 9058 8414 9534 8442
rect 9562 8414 9567 8442
rect 9646 8414 11382 8442
rect 11410 8414 11606 8442
rect 11634 8414 11639 8442
rect 12670 8414 13622 8442
rect 13650 8414 13846 8442
rect 13874 8414 13879 8442
rect 9646 8386 9674 8414
rect 12670 8386 12698 8414
rect 8969 8358 8974 8386
rect 9002 8358 9674 8386
rect 10649 8358 10654 8386
rect 10682 8358 11214 8386
rect 11242 8358 11247 8386
rect 12665 8358 12670 8386
rect 12698 8358 12703 8386
rect 12782 8358 13790 8386
rect 13818 8358 14574 8386
rect 14602 8358 14607 8386
rect 12782 8330 12810 8358
rect 9025 8302 9030 8330
rect 9058 8302 9422 8330
rect 9450 8302 10598 8330
rect 10626 8302 10631 8330
rect 11153 8302 11158 8330
rect 11186 8302 12782 8330
rect 12810 8302 12815 8330
rect 13225 8302 13230 8330
rect 13258 8302 13846 8330
rect 13874 8302 13879 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 0 8106 400 8120
rect 20600 8106 21000 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 6729 8078 6734 8106
rect 6762 8078 8526 8106
rect 8554 8078 8559 8106
rect 11489 8078 11494 8106
rect 11522 8078 12614 8106
rect 12642 8078 12647 8106
rect 20001 8078 20006 8106
rect 20034 8078 21000 8106
rect 0 8064 400 8078
rect 20600 8064 21000 8078
rect 8353 8022 8358 8050
rect 8386 8022 8414 8050
rect 8442 8022 8447 8050
rect 11881 8022 11886 8050
rect 11914 8022 12502 8050
rect 12530 8022 12726 8050
rect 12754 8022 13062 8050
rect 13090 8022 13095 8050
rect 12217 7910 12222 7938
rect 12250 7910 12726 7938
rect 12754 7910 13174 7938
rect 13202 7910 13207 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 12665 7798 12670 7826
rect 12698 7798 12703 7826
rect 12670 7770 12698 7798
rect 10313 7742 10318 7770
rect 10346 7742 10878 7770
rect 10906 7742 13062 7770
rect 13090 7742 13095 7770
rect 9081 7630 9086 7658
rect 9114 7630 9422 7658
rect 9450 7630 9455 7658
rect 8129 7574 8134 7602
rect 8162 7574 8974 7602
rect 9002 7574 9007 7602
rect 10985 7574 10990 7602
rect 11018 7574 11830 7602
rect 11858 7574 11863 7602
rect 11998 7546 12026 7742
rect 12497 7686 12502 7714
rect 12530 7686 12670 7714
rect 12698 7686 12703 7714
rect 13062 7658 13090 7742
rect 13062 7630 14294 7658
rect 14322 7630 14742 7658
rect 14770 7630 14775 7658
rect 13953 7574 13958 7602
rect 13986 7574 14518 7602
rect 14546 7574 18830 7602
rect 18858 7574 18863 7602
rect 11993 7518 11998 7546
rect 12026 7518 12031 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 9305 7294 9310 7322
rect 9338 7294 9478 7322
rect 9506 7294 10178 7322
rect 10150 7266 10178 7294
rect 7793 7238 7798 7266
rect 7826 7238 8246 7266
rect 8274 7238 9366 7266
rect 9394 7238 9702 7266
rect 9730 7238 9735 7266
rect 10145 7238 10150 7266
rect 10178 7238 13118 7266
rect 13146 7238 13151 7266
rect 8465 7182 8470 7210
rect 8498 7182 8974 7210
rect 9002 7182 10766 7210
rect 10794 7182 10799 7210
rect 9193 7126 9198 7154
rect 9226 7126 9422 7154
rect 9450 7126 9455 7154
rect 10089 7070 10094 7098
rect 10122 7070 10127 7098
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 10094 6986 10122 7070
rect 10033 6958 10038 6986
rect 10066 6958 10122 6986
rect 11993 6958 11998 6986
rect 12026 6958 12614 6986
rect 12642 6958 12647 6986
rect 10089 6846 10094 6874
rect 10122 6846 10127 6874
rect 8129 6790 8134 6818
rect 8162 6790 8862 6818
rect 8890 6790 8895 6818
rect 10094 6706 10122 6846
rect 13057 6790 13062 6818
rect 13090 6790 14070 6818
rect 14098 6790 14103 6818
rect 10094 6678 10878 6706
rect 10906 6678 10911 6706
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 9417 2030 9422 2058
rect 9450 2030 10038 2058
rect 10066 2030 10071 2058
rect 12105 2030 12110 2058
rect 12138 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 10761 1806 10766 1834
rect 10794 1806 11214 1834
rect 11242 1806 11247 1834
rect 11769 1806 11774 1834
rect 11802 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 8862 9758 8890 9786
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 8414 9310 8442 9338
rect 8862 9198 8890 9226
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 8414 8022 8442 8050
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 2224 9030 2384 9786
rect 8862 9786 8890 9791
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 8414 9338 8442 9343
rect 8414 8050 8442 9310
rect 8862 9226 8890 9758
rect 8862 9193 8890 9198
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 8414 8017 8442 8022
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7616 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7896 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _109_
timestamp 1698175906
transform 1 0 7168 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform -1 0 7672 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _111_
timestamp 1698175906
transform 1 0 11704 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8904 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform 1 0 8568 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10136 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11480 0 -1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11872 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 12880 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12824 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_
timestamp 1698175906
transform -1 0 10136 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _121_
timestamp 1698175906
transform -1 0 11032 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform -1 0 10920 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11928 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10640 0 -1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 12880 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1698175906
transform -1 0 10248 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _127_
timestamp 1698175906
transform 1 0 8904 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _128_
timestamp 1698175906
transform 1 0 10136 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698175906
transform -1 0 10472 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _130_
timestamp 1698175906
transform 1 0 10024 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _131_
timestamp 1698175906
transform 1 0 7952 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8792 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _134_
timestamp 1698175906
transform -1 0 9296 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _135_
timestamp 1698175906
transform -1 0 9576 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _136_
timestamp 1698175906
transform 1 0 7280 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform 1 0 8232 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 9240 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11032 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9632 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _141_
timestamp 1698175906
transform -1 0 9128 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _142_
timestamp 1698175906
transform 1 0 11032 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9520 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform 1 0 8176 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 13216 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _146_
timestamp 1698175906
transform 1 0 11032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 12936 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _148_
timestamp 1698175906
transform -1 0 12936 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7336 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _150_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7448 0 -1 10976
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _151_
timestamp 1698175906
transform -1 0 6328 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _152_
timestamp 1698175906
transform -1 0 9912 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _153_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10080 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 8624 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 12432 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform -1 0 12152 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_
timestamp 1698175906
transform 1 0 12208 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _158_
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13552 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _160_
timestamp 1698175906
transform -1 0 13608 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _161_
timestamp 1698175906
transform 1 0 10192 0 -1 11760
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _162_
timestamp 1698175906
transform 1 0 13104 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform -1 0 13888 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform -1 0 9408 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _165_
timestamp 1698175906
transform 1 0 8736 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _166_
timestamp 1698175906
transform -1 0 9352 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform 1 0 10024 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _168_
timestamp 1698175906
transform 1 0 12768 0 -1 13328
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _169_
timestamp 1698175906
transform -1 0 13048 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _170_
timestamp 1698175906
transform -1 0 11312 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _171_
timestamp 1698175906
transform 1 0 12880 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform 1 0 14112 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform -1 0 14112 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _174_
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _175_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14280 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _176_
timestamp 1698175906
transform -1 0 11872 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _177_
timestamp 1698175906
transform 1 0 12432 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _178_
timestamp 1698175906
transform 1 0 11144 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _179_
timestamp 1698175906
transform 1 0 11816 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _180_
timestamp 1698175906
transform -1 0 11032 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _181_
timestamp 1698175906
transform -1 0 8736 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9184 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _183_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10136 0 -1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _184_
timestamp 1698175906
transform -1 0 9632 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11088 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _186_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _187_
timestamp 1698175906
transform -1 0 9240 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _189_
timestamp 1698175906
transform 1 0 13720 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _190_
timestamp 1698175906
transform 1 0 12880 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11424 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform 1 0 7840 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _193_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7728 0 -1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _194_
timestamp 1698175906
transform -1 0 7672 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _195_
timestamp 1698175906
transform -1 0 8792 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698175906
transform -1 0 8904 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11368 0 1 9408
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _198_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9520 0 -1 10976
box -43 -43 2059 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _199_
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _200_
timestamp 1698175906
transform 1 0 8400 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _201_
timestamp 1698175906
transform -1 0 8568 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _202_
timestamp 1698175906
transform -1 0 7840 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _203_
timestamp 1698175906
transform 1 0 10192 0 1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _204_
timestamp 1698175906
transform -1 0 10248 0 -1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _205_
timestamp 1698175906
transform 1 0 9912 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _206_
timestamp 1698175906
transform 1 0 13160 0 -1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13440 0 1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _208_
timestamp 1698175906
transform 1 0 8120 0 -1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _209_
timestamp 1698175906
transform 1 0 7952 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _210_
timestamp 1698175906
transform -1 0 7784 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _211_
timestamp 1698175906
transform -1 0 10080 0 1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _212_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9800 0 1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _213_
timestamp 1698175906
transform 1 0 9464 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11144 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 9520 0 -1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 7672 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 5544 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 5376 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 6664 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform -1 0 12936 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 13608 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _223_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12936 0 -1 12544
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 7672 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 11984 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 14392 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 13720 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 10808 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 10248 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform -1 0 8288 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 10416 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 12992 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform -1 0 7448 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 6888 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform -1 0 8064 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 9520 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 12768 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 8848 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _242_
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _243_
timestamp 1698175906
transform 1 0 14056 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12768 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 9688 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 7000 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 12936 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 13496 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 14784 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 9408 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform -1 0 13720 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 14280 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 13608 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 11984 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform -1 0 12264 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 14728 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 7560 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform -1 0 9128 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 8176 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform -1 0 9520 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 14616 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 8288 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 11536 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11592 0 1 9408
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698175906
transform 1 0 9072 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698175906
transform 1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698175906
transform 1 0 9408 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_183 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10920 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_199
timestamp 1698175906
transform 1 0 11816 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_209
timestamp 1698175906
transform 1 0 12376 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698175906
transform 1 0 14280 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_150
timestamp 1698175906
transform 1 0 9072 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_154
timestamp 1698175906
transform 1 0 9296 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_187
timestamp 1698175906
transform 1 0 11144 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_203
timestamp 1698175906
transform 1 0 12040 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_207
timestamp 1698175906
transform 1 0 12264 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698175906
transform 1 0 12376 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_123
timestamp 1698175906
transform 1 0 7560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_154
timestamp 1698175906
transform 1 0 9296 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_158
timestamp 1698175906
transform 1 0 9520 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_152
timestamp 1698175906
transform 1 0 9184 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_160
timestamp 1698175906
transform 1 0 9632 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_164
timestamp 1698175906
transform 1 0 9856 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_200
timestamp 1698175906
transform 1 0 11872 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_204
timestamp 1698175906
transform 1 0 12096 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_208
timestamp 1698175906
transform 1 0 12320 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_241
timestamp 1698175906
transform 1 0 14168 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_245
timestamp 1698175906
transform 1 0 14392 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698175906
transform 1 0 16184 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 16296 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_159
timestamp 1698175906
transform 1 0 9576 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_163
timestamp 1698175906
transform 1 0 9800 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_185
timestamp 1698175906
transform 1 0 11032 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_201
timestamp 1698175906
transform 1 0 11928 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_209
timestamp 1698175906
transform 1 0 12376 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_224
timestamp 1698175906
transform 1 0 13216 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 14112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_156
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_188
timestamp 1698175906
transform 1 0 11200 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_196
timestamp 1698175906
transform 1 0 11648 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_198
timestamp 1698175906
transform 1 0 11760 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 12264 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_219
timestamp 1698175906
transform 1 0 12936 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_249
timestamp 1698175906
transform 1 0 14616 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_253
timestamp 1698175906
transform 1 0 14840 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_269
timestamp 1698175906
transform 1 0 15736 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698175906
transform 1 0 16184 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_144
timestamp 1698175906
transform 1 0 8736 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_160
timestamp 1698175906
transform 1 0 9632 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_168
timestamp 1698175906
transform 1 0 10080 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_224
timestamp 1698175906
transform 1 0 13216 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_232
timestamp 1698175906
transform 1 0 13664 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_239
timestamp 1698175906
transform 1 0 14056 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 14280 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_106
timestamp 1698175906
transform 1 0 6608 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_136
timestamp 1698175906
transform 1 0 8288 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_160
timestamp 1698175906
transform 1 0 9632 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_176
timestamp 1698175906
transform 1 0 10528 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_183
timestamp 1698175906
transform 1 0 10920 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_195
timestamp 1698175906
transform 1 0 11592 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_203
timestamp 1698175906
transform 1 0 12040 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_216
timestamp 1698175906
transform 1 0 12768 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_228
timestamp 1698175906
transform 1 0 13440 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_230
timestamp 1698175906
transform 1 0 13552 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_262
timestamp 1698175906
transform 1 0 15344 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 16240 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698175906
transform 1 0 7560 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_131
timestamp 1698175906
transform 1 0 8008 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_135
timestamp 1698175906
transform 1 0 8232 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_153
timestamp 1698175906
transform 1 0 9240 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_193
timestamp 1698175906
transform 1 0 11480 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_201
timestamp 1698175906
transform 1 0 11928 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_205
timestamp 1698175906
transform 1 0 12152 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_212
timestamp 1698175906
transform 1 0 12544 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_228
timestamp 1698175906
transform 1 0 13440 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_231
timestamp 1698175906
transform 1 0 13608 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698175906
transform 1 0 14280 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_253
timestamp 1698175906
transform 1 0 14840 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_285
timestamp 1698175906
transform 1 0 16632 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_301
timestamp 1698175906
transform 1 0 17528 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_309
timestamp 1698175906
transform 1 0 17976 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698175906
transform 1 0 18200 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698175906
transform 1 0 5376 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_86
timestamp 1698175906
transform 1 0 5488 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_116
timestamp 1698175906
transform 1 0 7168 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_120
timestamp 1698175906
transform 1 0 7392 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 8288 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_155
timestamp 1698175906
transform 1 0 9352 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_178
timestamp 1698175906
transform 1 0 10640 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_224
timestamp 1698175906
transform 1 0 13216 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_260
timestamp 1698175906
transform 1 0 15232 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 16128 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698175906
transform 1 0 6888 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_115
timestamp 1698175906
transform 1 0 7112 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_117
timestamp 1698175906
transform 1 0 7224 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_131
timestamp 1698175906
transform 1 0 8008 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_168
timestamp 1698175906
transform 1 0 10080 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_191
timestamp 1698175906
transform 1 0 11368 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 5152 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_113
timestamp 1698175906
transform 1 0 7000 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_115
timestamp 1698175906
transform 1 0 7112 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_158
timestamp 1698175906
transform 1 0 9520 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_192
timestamp 1698175906
transform 1 0 11424 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_196
timestamp 1698175906
transform 1 0 11648 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_218
timestamp 1698175906
transform 1 0 12880 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_222
timestamp 1698175906
transform 1 0 13104 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_238
timestamp 1698175906
transform 1 0 14000 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_270
timestamp 1698175906
transform 1 0 15792 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_85
timestamp 1698175906
transform 1 0 5432 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_93
timestamp 1698175906
transform 1 0 5880 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 6888 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_227
timestamp 1698175906
transform 1 0 13384 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_231
timestamp 1698175906
transform 1 0 13608 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_251
timestamp 1698175906
transform 1 0 14728 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_104
timestamp 1698175906
transform 1 0 6496 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_108
timestamp 1698175906
transform 1 0 6720 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_129
timestamp 1698175906
transform 1 0 7896 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_153
timestamp 1698175906
transform 1 0 9240 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_157
timestamp 1698175906
transform 1 0 9464 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_205
timestamp 1698175906
transform 1 0 12152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_274
timestamp 1698175906
transform 1 0 16016 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_115
timestamp 1698175906
transform 1 0 7112 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_125
timestamp 1698175906
transform 1 0 7672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_127
timestamp 1698175906
transform 1 0 7784 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_133
timestamp 1698175906
transform 1 0 8120 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_228
timestamp 1698175906
transform 1 0 13440 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_236
timestamp 1698175906
transform 1 0 13888 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_240
timestamp 1698175906
transform 1 0 14112 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_242
timestamp 1698175906
transform 1 0 14224 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 2240 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 4032 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 4480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_121
timestamp 1698175906
transform 1 0 7448 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_125
timestamp 1698175906
transform 1 0 7672 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698175906
transform 1 0 8848 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698175906
transform 1 0 8960 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_183
timestamp 1698175906
transform 1 0 10920 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_191
timestamp 1698175906
transform 1 0 11368 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_201
timestamp 1698175906
transform 1 0 11928 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_217
timestamp 1698175906
transform 1 0 12824 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_221
timestamp 1698175906
transform 1 0 13048 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_253
timestamp 1698175906
transform 1 0 14840 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_269
timestamp 1698175906
transform 1 0 15736 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698175906
transform 1 0 7112 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_119
timestamp 1698175906
transform 1 0 7336 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_121
timestamp 1698175906
transform 1 0 7448 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_128
timestamp 1698175906
transform 1 0 7840 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_141
timestamp 1698175906
transform 1 0 8568 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_149
timestamp 1698175906
transform 1 0 9016 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_163
timestamp 1698175906
transform 1 0 9800 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 10304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698175906
transform 1 0 11032 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_221
timestamp 1698175906
transform 1 0 13048 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_229
timestamp 1698175906
transform 1 0 13496 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_96
timestamp 1698175906
transform 1 0 6048 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_100
timestamp 1698175906
transform 1 0 6272 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_102
timestamp 1698175906
transform 1 0 6384 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_132
timestamp 1698175906
transform 1 0 8064 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_149
timestamp 1698175906
transform 1 0 9016 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_157
timestamp 1698175906
transform 1 0 9464 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698175906
transform 1 0 9688 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_163
timestamp 1698175906
transform 1 0 9800 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_171
timestamp 1698175906
transform 1 0 10248 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_203
timestamp 1698175906
transform 1 0 12040 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698175906
transform 1 0 12264 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_218
timestamp 1698175906
transform 1 0 12880 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_250
timestamp 1698175906
transform 1 0 14672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_254
timestamp 1698175906
transform 1 0 14896 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_270
timestamp 1698175906
transform 1 0 15792 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_131
timestamp 1698175906
transform 1 0 8008 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_135
timestamp 1698175906
transform 1 0 8232 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_138
timestamp 1698175906
transform 1 0 8400 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_145
timestamp 1698175906
transform 1 0 8792 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_161
timestamp 1698175906
transform 1 0 9688 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_169
timestamp 1698175906
transform 1 0 10136 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698175906
transform 1 0 10360 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_186
timestamp 1698175906
transform 1 0 11088 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_236
timestamp 1698175906
transform 1 0 13888 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_238
timestamp 1698175906
transform 1 0 14000 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_253
timestamp 1698175906
transform 1 0 14840 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_285
timestamp 1698175906
transform 1 0 16632 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_301
timestamp 1698175906
transform 1 0 17528 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698175906
transform 1 0 17976 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698175906
transform 1 0 18200 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_120
timestamp 1698175906
transform 1 0 7392 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_127
timestamp 1698175906
transform 1 0 7784 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_129
timestamp 1698175906
transform 1 0 7896 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 8400 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_146
timestamp 1698175906
transform 1 0 8848 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_153
timestamp 1698175906
transform 1 0 9240 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_173
timestamp 1698175906
transform 1 0 10360 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_203
timestamp 1698175906
transform 1 0 12040 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 12264 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_223
timestamp 1698175906
transform 1 0 13160 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_233
timestamp 1698175906
transform 1 0 13720 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_265
timestamp 1698175906
transform 1 0 15512 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 15960 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_136
timestamp 1698175906
transform 1 0 8288 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_183
timestamp 1698175906
transform 1 0 10920 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_215
timestamp 1698175906
transform 1 0 12712 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_231
timestamp 1698175906
transform 1 0 13608 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698175906
transform 1 0 14056 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 14280 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_108
timestamp 1698175906
transform 1 0 6720 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_110
timestamp 1698175906
transform 1 0 6832 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_147
timestamp 1698175906
transform 1 0 8904 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_151
timestamp 1698175906
transform 1 0 9128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_155
timestamp 1698175906
transform 1 0 9352 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_187
timestamp 1698175906
transform 1 0 11144 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_203
timestamp 1698175906
transform 1 0 12040 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 12264 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_139
timestamp 1698175906
transform 1 0 8456 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_155
timestamp 1698175906
transform 1 0 9352 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_168
timestamp 1698175906
transform 1 0 10080 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_168
timestamp 1698175906
transform 1 0 10080 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_195
timestamp 1698175906
transform 1 0 11592 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_203
timestamp 1698175906
transform 1 0 12040 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_40
timestamp 1698175906
transform 1 0 2912 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_42
timestamp 1698175906
transform 1 0 3024 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_47
timestamp 1698175906
transform 1 0 3304 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_63
timestamp 1698175906
transform 1 0 4200 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_67
timestamp 1698175906
transform 1 0 4424 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita42_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 3304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita42_26
timestamp 1698175906
transform -1 0 10640 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 10136 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 2240 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform -1 0 14280 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 9464 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 10640 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 3024 20600 3080 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 8064 20600 8120 21000 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 10080 20600 10136 21000 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 12096 0 12152 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 11424 400 11480 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 12768 0 12824 400 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 9408 0 9464 400 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 10752 0 10808 400 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 13020 6944 13020 6944 0 _000_
rlabel metal2 7084 10248 7084 10248 0 _001_
rlabel metal2 5964 10276 5964 10276 0 _002_
rlabel metal2 7140 8596 7140 8596 0 _003_
rlabel metal2 11984 10668 11984 10668 0 _004_
rlabel metal3 13776 9156 13776 9156 0 _005_
rlabel metal2 13412 12516 13412 12516 0 _006_
rlabel metal2 8148 6664 8148 6664 0 _007_
rlabel metal2 12796 12012 12796 12012 0 _008_
rlabel metal2 13972 10584 13972 10584 0 _009_
rlabel metal2 14168 8484 14168 8484 0 _010_
rlabel metal2 11284 8232 11284 8232 0 _011_
rlabel metal2 10724 6944 10724 6944 0 _012_
rlabel metal2 7812 8316 7812 8316 0 _013_
rlabel metal2 10864 13580 10864 13580 0 _014_
rlabel metal2 13356 8120 13356 8120 0 _015_
rlabel metal2 7420 11312 7420 11312 0 _016_
rlabel metal2 8540 13720 8540 13720 0 _017_
rlabel metal2 7588 12180 7588 12180 0 _018_
rlabel metal2 10080 13244 10080 13244 0 _019_
rlabel metal2 13216 10836 13216 10836 0 _020_
rlabel metal2 7140 13412 7140 13412 0 _021_
rlabel metal2 9464 13468 9464 13468 0 _022_
rlabel metal2 11760 11676 11760 11676 0 _023_
rlabel metal2 9996 6160 9996 6160 0 _024_
rlabel metal3 8568 7588 8568 7588 0 _025_
rlabel metal2 12180 10444 12180 10444 0 _026_
rlabel metal2 13356 9072 13356 9072 0 _027_
rlabel metal2 13860 9996 13860 9996 0 _028_
rlabel metal2 13524 9464 13524 9464 0 _029_
rlabel metal2 13748 12376 13748 12376 0 _030_
rlabel metal2 13356 12348 13356 12348 0 _031_
rlabel metal2 9044 6748 9044 6748 0 _032_
rlabel metal2 10220 11956 10220 11956 0 _033_
rlabel metal3 11592 11844 11592 11844 0 _034_
rlabel metal2 12964 12488 12964 12488 0 _035_
rlabel metal2 13860 10780 13860 10780 0 _036_
rlabel metal3 12488 7924 12488 7924 0 _037_
rlabel metal2 14168 10500 14168 10500 0 _038_
rlabel metal3 14420 8820 14420 8820 0 _039_
rlabel metal3 10528 8428 10528 8428 0 _040_
rlabel metal2 12600 8036 12600 8036 0 _041_
rlabel metal3 11424 7588 11424 7588 0 _042_
rlabel metal2 8652 7924 8652 7924 0 _043_
rlabel metal2 9548 11172 9548 11172 0 _044_
rlabel metal3 9800 12628 9800 12628 0 _045_
rlabel metal2 10780 13104 10780 13104 0 _046_
rlabel metal2 7532 11396 7532 11396 0 _047_
rlabel metal2 8764 13454 8764 13454 0 _048_
rlabel metal2 13860 8204 13860 8204 0 _049_
rlabel metal2 10780 10332 10780 10332 0 _050_
rlabel metal2 8008 11284 8008 11284 0 _051_
rlabel metal2 7616 11284 7616 11284 0 _052_
rlabel metal2 8820 14084 8820 14084 0 _053_
rlabel metal2 8652 13720 8652 13720 0 _054_
rlabel metal2 11172 10248 11172 10248 0 _055_
rlabel metal3 9660 11900 9660 11900 0 _056_
rlabel metal2 8624 12516 8624 12516 0 _057_
rlabel metal2 8204 11984 8204 11984 0 _058_
rlabel metal2 10304 13468 10304 13468 0 _059_
rlabel metal2 9940 12908 9940 12908 0 _060_
rlabel metal2 13300 10556 13300 10556 0 _061_
rlabel metal2 8344 13132 8344 13132 0 _062_
rlabel metal2 7896 13020 7896 13020 0 _063_
rlabel metal2 9772 14196 9772 14196 0 _064_
rlabel metal2 9548 12572 9548 12572 0 _065_
rlabel metal2 9268 9996 9268 9996 0 _066_
rlabel metal3 11508 11116 11508 11116 0 _067_
rlabel metal2 7532 10164 7532 10164 0 _068_
rlabel metal2 7420 10192 7420 10192 0 _069_
rlabel metal2 10948 9436 10948 9436 0 _070_
rlabel metal3 9156 9268 9156 9268 0 _071_
rlabel metal2 10276 9268 10276 9268 0 _072_
rlabel metal2 10276 8904 10276 8904 0 _073_
rlabel metal3 11928 10836 11928 10836 0 _074_
rlabel metal2 13020 8624 13020 8624 0 _075_
rlabel metal2 13300 12236 13300 12236 0 _076_
rlabel metal3 12236 11564 12236 11564 0 _077_
rlabel metal2 10780 9016 10780 9016 0 _078_
rlabel metal2 10976 9156 10976 9156 0 _079_
rlabel metal2 10836 9044 10836 9044 0 _080_
rlabel metal2 10836 11592 10836 11592 0 _081_
rlabel metal2 9884 11396 9884 11396 0 _082_
rlabel metal2 10164 7084 10164 7084 0 _083_
rlabel metal2 9996 6944 9996 6944 0 _084_
rlabel metal2 9940 11536 9940 11536 0 _085_
rlabel metal2 10360 8148 10360 8148 0 _086_
rlabel metal2 10360 7924 10360 7924 0 _087_
rlabel metal2 8988 10388 8988 10388 0 _088_
rlabel metal3 9380 11172 9380 11172 0 _089_
rlabel metal2 10108 11732 10108 11732 0 _090_
rlabel metal2 9044 10724 9044 10724 0 _091_
rlabel metal3 9268 7644 9268 7644 0 _092_
rlabel metal2 8372 9548 8372 9548 0 _093_
rlabel metal2 12348 9632 12348 9632 0 _094_
rlabel metal2 8988 8624 8988 8624 0 _095_
rlabel metal2 13972 8708 13972 8708 0 _096_
rlabel metal2 8820 8456 8820 8456 0 _097_
rlabel metal2 13468 9520 13468 9520 0 _098_
rlabel metal3 8484 9996 8484 9996 0 _099_
rlabel metal2 12964 11116 12964 11116 0 _100_
rlabel metal2 12908 7196 12908 7196 0 _101_
rlabel metal2 13804 8260 13804 8260 0 _102_
rlabel metal3 12796 8036 12796 8036 0 _103_
rlabel metal2 6244 10556 6244 10556 0 _104_
rlabel metal2 9940 9632 9940 9632 0 _105_
rlabel metal2 8568 8820 8568 8820 0 _106_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal2 11844 9968 11844 9968 0 clknet_0_clk
rlabel metal2 7364 11536 7364 11536 0 clknet_1_0__leaf_clk
rlabel metal2 13692 12824 13692 12824 0 clknet_1_1__leaf_clk
rlabel metal2 7084 9324 7084 9324 0 dut42.count\[0\]
rlabel metal2 7336 9996 7336 9996 0 dut42.count\[1\]
rlabel metal3 9128 8820 9128 8820 0 dut42.count\[2\]
rlabel metal3 11592 10052 11592 10052 0 dut42.count\[3\]
rlabel metal2 6748 8260 6748 8260 0 net1
rlabel metal2 8428 13944 8428 13944 0 net10
rlabel metal2 6524 12516 6524 12516 0 net11
rlabel metal2 11060 14056 11060 14056 0 net12
rlabel metal2 15260 8596 15260 8596 0 net13
rlabel metal2 12124 15960 12124 15960 0 net14
rlabel metal2 13972 7812 13972 7812 0 net15
rlabel metal2 15932 10556 15932 10556 0 net16
rlabel metal3 14742 12796 14742 12796 0 net17
rlabel metal2 9212 4144 9212 4144 0 net18
rlabel metal2 15148 9576 15148 9576 0 net19
rlabel metal2 14308 10696 14308 10696 0 net2
rlabel metal2 13972 3374 13972 3374 0 net20
rlabel metal2 9436 7056 9436 7056 0 net21
rlabel metal3 15960 11984 15960 11984 0 net22
rlabel metal2 11060 5964 11060 5964 0 net23
rlabel metal2 18956 12908 18956 12908 0 net24
rlabel metal2 3108 18956 3108 18956 0 net25
rlabel metal2 10472 18956 10472 18956 0 net26
rlabel metal2 8204 13888 8204 13888 0 net3
rlabel metal2 10388 13888 10388 13888 0 net4
rlabel metal2 18788 13076 18788 13076 0 net5
rlabel metal2 12040 7644 12040 7644 0 net6
rlabel metal2 12348 7952 12348 7952 0 net7
rlabel metal2 14588 12460 14588 12460 0 net8
rlabel metal2 5908 11536 5908 11536 0 net9
rlabel metal3 679 8092 679 8092 0 segm[10]
rlabel metal2 20020 11004 20020 11004 0 segm[11]
rlabel metal2 8092 19677 8092 19677 0 segm[12]
rlabel metal2 10108 19677 10108 19677 0 segm[13]
rlabel metal2 20020 13356 20020 13356 0 segm[1]
rlabel metal3 12292 1820 12292 1820 0 segm[2]
rlabel metal3 12628 2044 12628 2044 0 segm[3]
rlabel metal2 20020 12180 20020 12180 0 segm[5]
rlabel metal3 679 11452 679 11452 0 segm[6]
rlabel metal2 8764 19873 8764 19873 0 segm[7]
rlabel metal3 679 12460 679 12460 0 segm[8]
rlabel metal2 10780 19873 10780 19873 0 segm[9]
rlabel metal2 20020 8820 20020 8820 0 sel[0]
rlabel metal2 11788 19873 11788 19873 0 sel[10]
rlabel metal2 20020 8204 20020 8204 0 sel[11]
rlabel metal2 20020 10556 20020 10556 0 sel[1]
rlabel metal2 20020 12628 20020 12628 0 sel[2]
rlabel metal2 9100 1029 9100 1029 0 sel[3]
rlabel metal2 20020 9548 20020 9548 0 sel[4]
rlabel metal2 12796 427 12796 427 0 sel[5]
rlabel metal3 9744 2044 9744 2044 0 sel[6]
rlabel metal2 20020 11900 20020 11900 0 sel[7]
rlabel metal3 11004 1820 11004 1820 0 sel[8]
rlabel metal2 19964 12936 19964 12936 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
