magic
tech gf180mcuD
magscale 1 5
timestamp 1699641524
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9031 19137 9057 19143
rect 9031 19105 9057 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 8521 18999 8527 19025
rect 8553 18999 8559 19025
rect 10873 18999 10879 19025
rect 10905 18999 10911 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 9983 18969 10009 18975
rect 9983 18937 10009 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 10039 18745 10065 18751
rect 10039 18713 10065 18719
rect 13735 18745 13761 18751
rect 13735 18713 13761 18719
rect 9529 18607 9535 18633
rect 9561 18607 9567 18633
rect 13393 18607 13399 18633
rect 13425 18607 13431 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 20119 18129 20145 18135
rect 20119 18097 20145 18103
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 11663 14041 11689 14047
rect 11663 14009 11689 14015
rect 11551 13929 11577 13935
rect 11551 13897 11577 13903
rect 11719 13929 11745 13935
rect 11719 13897 11745 13903
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 9529 13567 9535 13593
rect 9561 13567 9567 13593
rect 12105 13567 12111 13593
rect 12137 13567 12143 13593
rect 9815 13537 9841 13543
rect 8073 13511 8079 13537
rect 8105 13511 8111 13537
rect 10705 13511 10711 13537
rect 10737 13511 10743 13537
rect 9815 13505 9841 13511
rect 9647 13481 9673 13487
rect 8465 13455 8471 13481
rect 8497 13455 8503 13481
rect 9647 13449 9673 13455
rect 9759 13481 9785 13487
rect 11041 13455 11047 13481
rect 11073 13455 11079 13481
rect 9759 13449 9785 13455
rect 12335 13425 12361 13431
rect 12335 13393 12361 13399
rect 20119 13425 20145 13431
rect 20119 13393 20145 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8695 13257 8721 13263
rect 8695 13225 8721 13231
rect 8807 13257 8833 13263
rect 8807 13225 8833 13231
rect 11551 13257 11577 13263
rect 11551 13225 11577 13231
rect 11831 13201 11857 13207
rect 11831 13169 11857 13175
rect 8863 13145 8889 13151
rect 11495 13145 11521 13151
rect 11265 13119 11271 13145
rect 11297 13119 11303 13145
rect 8863 13113 8889 13119
rect 11495 13113 11521 13119
rect 12671 13089 12697 13095
rect 9865 13063 9871 13089
rect 9897 13063 9903 13089
rect 10929 13063 10935 13089
rect 10961 13063 10967 13089
rect 12671 13057 12697 13063
rect 11551 13033 11577 13039
rect 11551 13001 11577 13007
rect 12615 13033 12641 13039
rect 12615 13001 12641 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 10935 12865 10961 12871
rect 10935 12833 10961 12839
rect 8353 12783 8359 12809
rect 8385 12783 8391 12809
rect 12329 12783 12335 12809
rect 12361 12783 12367 12809
rect 13393 12783 13399 12809
rect 13425 12783 13431 12809
rect 6953 12727 6959 12753
rect 6985 12727 6991 12753
rect 11937 12727 11943 12753
rect 11969 12727 11975 12753
rect 8583 12697 8609 12703
rect 7289 12671 7295 12697
rect 7321 12671 7327 12697
rect 8583 12665 8609 12671
rect 8639 12697 8665 12703
rect 8639 12665 8665 12671
rect 9031 12697 9057 12703
rect 10655 12697 10681 12703
rect 9193 12671 9199 12697
rect 9225 12671 9231 12697
rect 9031 12665 9057 12671
rect 10655 12665 10681 12671
rect 10879 12697 10905 12703
rect 10879 12665 10905 12671
rect 10991 12697 11017 12703
rect 10991 12665 11017 12671
rect 11103 12697 11129 12703
rect 11103 12665 11129 12671
rect 11159 12697 11185 12703
rect 11159 12665 11185 12671
rect 8471 12641 8497 12647
rect 8471 12609 8497 12615
rect 10767 12641 10793 12647
rect 10767 12609 10793 12615
rect 13623 12641 13649 12647
rect 13623 12609 13649 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 8135 12473 8161 12479
rect 8135 12441 8161 12447
rect 12167 12473 12193 12479
rect 12167 12441 12193 12447
rect 12223 12473 12249 12479
rect 12223 12441 12249 12447
rect 12279 12473 12305 12479
rect 12279 12441 12305 12447
rect 7967 12361 7993 12367
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 7065 12335 7071 12361
rect 7097 12335 7103 12361
rect 7967 12329 7993 12335
rect 8135 12361 8161 12367
rect 8135 12329 8161 12335
rect 8303 12361 8329 12367
rect 12111 12361 12137 12367
rect 9025 12335 9031 12361
rect 9057 12335 9063 12361
rect 11993 12335 11999 12361
rect 12025 12335 12031 12361
rect 8303 12329 8329 12335
rect 12111 12329 12137 12335
rect 5665 12279 5671 12305
rect 5697 12279 5703 12305
rect 6729 12279 6735 12305
rect 6761 12279 6767 12305
rect 9361 12279 9367 12305
rect 9393 12279 9399 12305
rect 10425 12279 10431 12305
rect 10457 12279 10463 12305
rect 967 12249 993 12255
rect 967 12217 993 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 7519 12025 7545 12031
rect 7519 11993 7545 11999
rect 9647 12025 9673 12031
rect 12951 12025 12977 12031
rect 12721 11999 12727 12025
rect 12753 11999 12759 12025
rect 9647 11993 9673 11999
rect 12951 11993 12977 11999
rect 20007 12025 20033 12031
rect 20007 11993 20033 11999
rect 7071 11969 7097 11975
rect 7071 11937 7097 11943
rect 7463 11969 7489 11975
rect 7625 11943 7631 11969
rect 7657 11943 7663 11969
rect 11265 11943 11271 11969
rect 11297 11943 11303 11969
rect 18937 11943 18943 11969
rect 18969 11943 18975 11969
rect 7463 11937 7489 11943
rect 13567 11913 13593 11919
rect 11657 11887 11663 11913
rect 11689 11887 11695 11913
rect 13567 11881 13593 11887
rect 7015 11857 7041 11863
rect 7015 11825 7041 11831
rect 7127 11857 7153 11863
rect 7127 11825 7153 11831
rect 7239 11857 7265 11863
rect 7239 11825 7265 11831
rect 9479 11857 9505 11863
rect 9479 11825 9505 11831
rect 9591 11857 9617 11863
rect 9591 11825 9617 11831
rect 9703 11857 9729 11863
rect 9703 11825 9729 11831
rect 13623 11857 13649 11863
rect 13623 11825 13649 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 10879 11689 10905 11695
rect 10879 11657 10905 11663
rect 11159 11689 11185 11695
rect 11159 11657 11185 11663
rect 11719 11689 11745 11695
rect 11719 11657 11745 11663
rect 12727 11689 12753 11695
rect 12727 11657 12753 11663
rect 8807 11633 8833 11639
rect 8807 11601 8833 11607
rect 8919 11633 8945 11639
rect 8919 11601 8945 11607
rect 9199 11633 9225 11639
rect 12671 11633 12697 11639
rect 10481 11607 10487 11633
rect 10513 11607 10519 11633
rect 9199 11601 9225 11607
rect 12671 11601 12697 11607
rect 12951 11633 12977 11639
rect 13673 11607 13679 11633
rect 13705 11607 13711 11633
rect 12951 11601 12977 11607
rect 9255 11577 9281 11583
rect 6953 11551 6959 11577
rect 6985 11551 6991 11577
rect 9255 11545 9281 11551
rect 9927 11577 9953 11583
rect 9927 11545 9953 11551
rect 10319 11577 10345 11583
rect 10319 11545 10345 11551
rect 10599 11577 10625 11583
rect 10761 11551 10767 11577
rect 10793 11551 10799 11577
rect 11041 11551 11047 11577
rect 11073 11551 11079 11577
rect 12777 11551 12783 11577
rect 12809 11551 12815 11577
rect 13337 11551 13343 11577
rect 13369 11551 13375 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 10599 11545 10625 11551
rect 8863 11521 8889 11527
rect 14967 11521 14993 11527
rect 7345 11495 7351 11521
rect 7377 11495 7383 11521
rect 8409 11495 8415 11521
rect 8441 11495 8447 11521
rect 10817 11495 10823 11521
rect 10849 11495 10855 11521
rect 11657 11495 11663 11521
rect 11689 11495 11695 11521
rect 14737 11495 14743 11521
rect 14769 11495 14775 11521
rect 8863 11489 8889 11495
rect 14967 11489 14993 11495
rect 9199 11465 9225 11471
rect 9199 11433 9225 11439
rect 9871 11465 9897 11471
rect 9871 11433 9897 11439
rect 11215 11465 11241 11471
rect 11215 11433 11241 11439
rect 11831 11465 11857 11471
rect 11831 11433 11857 11439
rect 13063 11465 13089 11471
rect 13063 11433 13089 11439
rect 13119 11465 13145 11471
rect 13119 11433 13145 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 967 11241 993 11247
rect 967 11209 993 11215
rect 8191 11241 8217 11247
rect 8191 11209 8217 11215
rect 11887 11241 11913 11247
rect 11887 11209 11913 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 6847 11185 6873 11191
rect 2137 11159 2143 11185
rect 2169 11159 2175 11185
rect 6847 11153 6873 11159
rect 6959 11185 6985 11191
rect 6959 11153 6985 11159
rect 7183 11185 7209 11191
rect 7183 11153 7209 11159
rect 8303 11185 8329 11191
rect 8303 11153 8329 11159
rect 8359 11185 8385 11191
rect 11495 11185 11521 11191
rect 10033 11159 10039 11185
rect 10065 11159 10071 11185
rect 10257 11159 10263 11185
rect 10289 11159 10295 11185
rect 11209 11159 11215 11185
rect 11241 11159 11247 11185
rect 8359 11153 8385 11159
rect 11495 11153 11521 11159
rect 11775 11185 11801 11191
rect 11775 11153 11801 11159
rect 11999 11185 12025 11191
rect 13623 11185 13649 11191
rect 12273 11159 12279 11185
rect 12305 11159 12311 11185
rect 13169 11159 13175 11185
rect 13201 11159 13207 11185
rect 13337 11159 13343 11185
rect 13369 11159 13375 11185
rect 11999 11153 12025 11159
rect 13623 11153 13649 11159
rect 13679 11185 13705 11191
rect 13679 11153 13705 11159
rect 14239 11185 14265 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 14239 11153 14265 11159
rect 8135 11129 8161 11135
rect 8135 11097 8161 11103
rect 9143 11129 9169 11135
rect 13455 11129 13481 11135
rect 9305 11103 9311 11129
rect 9337 11103 9343 11129
rect 9753 11103 9759 11129
rect 9785 11103 9791 11129
rect 9865 11103 9871 11129
rect 9897 11103 9903 11129
rect 10369 11103 10375 11129
rect 10401 11103 10407 11129
rect 11657 11103 11663 11129
rect 11689 11103 11695 11129
rect 9143 11097 9169 11103
rect 13455 11097 13481 11103
rect 14295 11129 14321 11135
rect 14295 11097 14321 11103
rect 6903 11073 6929 11079
rect 6903 11041 6929 11047
rect 8807 11073 8833 11079
rect 10711 11073 10737 11079
rect 11775 11073 11801 11079
rect 13287 11073 13313 11079
rect 8969 11047 8975 11073
rect 9001 11047 9007 11073
rect 9529 11047 9535 11073
rect 9561 11047 9567 11073
rect 10873 11047 10879 11073
rect 10905 11047 10911 11073
rect 11097 11047 11103 11073
rect 11129 11047 11135 11073
rect 12161 11047 12167 11073
rect 12193 11047 12199 11073
rect 8807 11041 8833 11047
rect 10711 11041 10737 11047
rect 11775 11041 11801 11047
rect 13287 11041 13313 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8807 10905 8833 10911
rect 9305 10879 9311 10905
rect 9337 10879 9343 10905
rect 8807 10873 8833 10879
rect 8359 10849 8385 10855
rect 8969 10823 8975 10849
rect 9001 10823 9007 10849
rect 8359 10817 8385 10823
rect 7071 10793 7097 10799
rect 6897 10767 6903 10793
rect 6929 10767 6935 10793
rect 7071 10761 7097 10767
rect 7239 10793 7265 10799
rect 7239 10761 7265 10767
rect 7407 10793 7433 10799
rect 9535 10793 9561 10799
rect 9193 10767 9199 10793
rect 9225 10767 9231 10793
rect 9753 10767 9759 10793
rect 9785 10767 9791 10793
rect 12609 10767 12615 10793
rect 12641 10767 12647 10793
rect 7407 10761 7433 10767
rect 9535 10761 9561 10767
rect 7295 10737 7321 10743
rect 5441 10711 5447 10737
rect 5473 10711 5479 10737
rect 6505 10711 6511 10737
rect 6537 10711 6543 10737
rect 11713 10711 11719 10737
rect 11745 10711 11751 10737
rect 15017 10711 15023 10737
rect 15049 10711 15055 10737
rect 7295 10705 7321 10711
rect 8415 10681 8441 10687
rect 8415 10649 8441 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 6735 10513 6761 10519
rect 6735 10481 6761 10487
rect 6903 10513 6929 10519
rect 6903 10481 6929 10487
rect 967 10457 993 10463
rect 12615 10457 12641 10463
rect 4993 10431 4999 10457
rect 5025 10431 5031 10457
rect 9025 10431 9031 10457
rect 9057 10431 9063 10457
rect 11769 10431 11775 10457
rect 11801 10431 11807 10457
rect 967 10425 993 10431
rect 12615 10425 12641 10431
rect 20007 10457 20033 10463
rect 20007 10425 20033 10431
rect 12391 10401 12417 10407
rect 2137 10375 2143 10401
rect 2169 10375 2175 10401
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 10761 10375 10767 10401
rect 10793 10375 10799 10401
rect 10929 10375 10935 10401
rect 10961 10375 10967 10401
rect 11377 10375 11383 10401
rect 11409 10375 11415 10401
rect 11881 10375 11887 10401
rect 11913 10375 11919 10401
rect 12391 10369 12417 10375
rect 12839 10401 12865 10407
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 12839 10369 12865 10375
rect 6791 10345 6817 10351
rect 12503 10345 12529 10351
rect 6057 10319 6063 10345
rect 6089 10319 6095 10345
rect 11153 10319 11159 10345
rect 11185 10319 11191 10345
rect 11433 10319 11439 10345
rect 11465 10319 11471 10345
rect 12161 10319 12167 10345
rect 12193 10319 12199 10345
rect 6791 10313 6817 10319
rect 12503 10313 12529 10319
rect 12671 10345 12697 10351
rect 13511 10345 13537 10351
rect 13001 10319 13007 10345
rect 13033 10319 13039 10345
rect 12671 10313 12697 10319
rect 13511 10313 13537 10319
rect 13567 10345 13593 10351
rect 13567 10313 13593 10319
rect 13679 10289 13705 10295
rect 10705 10263 10711 10289
rect 10737 10263 10743 10289
rect 13679 10257 13705 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 10263 10121 10289 10127
rect 10263 10089 10289 10095
rect 10991 10121 11017 10127
rect 10991 10089 11017 10095
rect 11103 10121 11129 10127
rect 11103 10089 11129 10095
rect 11943 10121 11969 10127
rect 11943 10089 11969 10095
rect 12727 10093 12753 10099
rect 6567 10065 6593 10071
rect 6567 10033 6593 10039
rect 6679 10065 6705 10071
rect 6679 10033 6705 10039
rect 6847 10065 6873 10071
rect 6847 10033 6873 10039
rect 6903 10065 6929 10071
rect 6903 10033 6929 10039
rect 9087 10065 9113 10071
rect 9087 10033 9113 10039
rect 10375 10065 10401 10071
rect 10375 10033 10401 10039
rect 11159 10065 11185 10071
rect 11159 10033 11185 10039
rect 11887 10065 11913 10071
rect 11887 10033 11913 10039
rect 11999 10065 12025 10071
rect 11999 10033 12025 10039
rect 12671 10065 12697 10071
rect 12727 10061 12753 10067
rect 12895 10065 12921 10071
rect 12671 10033 12697 10039
rect 13729 10039 13735 10065
rect 13761 10039 13767 10065
rect 12895 10033 12921 10039
rect 6511 10009 6537 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 6511 9977 6537 9983
rect 9423 10009 9449 10015
rect 10319 10009 10345 10015
rect 9585 9983 9591 10009
rect 9617 9983 9623 10009
rect 9423 9977 9449 9983
rect 10319 9977 10345 9983
rect 13007 10009 13033 10015
rect 13007 9977 13033 9983
rect 13231 10009 13257 10015
rect 13337 9983 13343 10009
rect 13369 9983 13375 10009
rect 13231 9977 13257 9983
rect 13119 9953 13145 9959
rect 15023 9953 15049 9959
rect 9137 9927 9143 9953
rect 9169 9927 9175 9953
rect 9865 9927 9871 9953
rect 9897 9927 9903 9953
rect 14793 9927 14799 9953
rect 14825 9927 14831 9953
rect 13119 9921 13145 9927
rect 15023 9921 15049 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 6847 9897 6873 9903
rect 6847 9865 6873 9871
rect 8975 9897 9001 9903
rect 12671 9897 12697 9903
rect 9529 9871 9535 9897
rect 9561 9871 9567 9897
rect 8975 9865 9001 9871
rect 12671 9865 12697 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 11215 9729 11241 9735
rect 11215 9697 11241 9703
rect 11943 9729 11969 9735
rect 11943 9697 11969 9703
rect 967 9673 993 9679
rect 4993 9647 4999 9673
rect 5025 9647 5031 9673
rect 9361 9647 9367 9673
rect 9393 9647 9399 9673
rect 13225 9647 13231 9673
rect 13257 9647 13263 9673
rect 14289 9647 14295 9673
rect 14321 9647 14327 9673
rect 967 9641 993 9647
rect 8807 9617 8833 9623
rect 10039 9617 10065 9623
rect 14575 9617 14601 9623
rect 2137 9591 2143 9617
rect 2169 9591 2175 9617
rect 6449 9591 6455 9617
rect 6481 9591 6487 9617
rect 9417 9591 9423 9617
rect 9449 9591 9455 9617
rect 9585 9591 9591 9617
rect 9617 9591 9623 9617
rect 11657 9591 11663 9617
rect 11689 9591 11695 9617
rect 12889 9591 12895 9617
rect 12921 9591 12927 9617
rect 8807 9585 8833 9591
rect 10039 9585 10065 9591
rect 14575 9585 14601 9591
rect 14687 9617 14713 9623
rect 14687 9585 14713 9591
rect 6903 9561 6929 9567
rect 6057 9535 6063 9561
rect 6089 9535 6095 9561
rect 6903 9529 6929 9535
rect 7071 9561 7097 9567
rect 11271 9561 11297 9567
rect 9193 9535 9199 9561
rect 9225 9535 9231 9561
rect 7071 9529 7097 9535
rect 11271 9529 11297 9535
rect 11775 9505 11801 9511
rect 8969 9479 8975 9505
rect 9001 9479 9007 9505
rect 9865 9479 9871 9505
rect 9897 9479 9903 9505
rect 11775 9473 11801 9479
rect 11887 9505 11913 9511
rect 11887 9473 11913 9479
rect 14631 9505 14657 9511
rect 14631 9473 14657 9479
rect 14799 9505 14825 9511
rect 14799 9473 14825 9479
rect 15079 9505 15105 9511
rect 15079 9473 15105 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 5895 9337 5921 9343
rect 9815 9337 9841 9343
rect 6505 9311 6511 9337
rect 6537 9311 6543 9337
rect 5895 9305 5921 9311
rect 9815 9305 9841 9311
rect 6399 9281 6425 9287
rect 6399 9249 6425 9255
rect 7127 9281 7153 9287
rect 7127 9249 7153 9255
rect 9759 9281 9785 9287
rect 9759 9249 9785 9255
rect 10151 9281 10177 9287
rect 10151 9249 10177 9255
rect 10879 9281 10905 9287
rect 10879 9249 10905 9255
rect 10935 9281 10961 9287
rect 11545 9255 11551 9281
rect 11577 9255 11583 9281
rect 10935 9249 10961 9255
rect 5839 9225 5865 9231
rect 5839 9193 5865 9199
rect 6567 9225 6593 9231
rect 7295 9225 7321 9231
rect 6785 9199 6791 9225
rect 6817 9199 6823 9225
rect 6567 9193 6593 9199
rect 7295 9193 7321 9199
rect 9255 9225 9281 9231
rect 9647 9225 9673 9231
rect 9417 9199 9423 9225
rect 9449 9199 9455 9225
rect 9255 9193 9281 9199
rect 9647 9193 9673 9199
rect 10039 9225 10065 9231
rect 10375 9225 10401 9231
rect 10313 9199 10319 9225
rect 10345 9199 10351 9225
rect 10039 9193 10065 9199
rect 10375 9193 10401 9199
rect 10431 9225 10457 9231
rect 10431 9193 10457 9199
rect 10767 9225 10793 9231
rect 11321 9199 11327 9225
rect 11353 9199 11359 9225
rect 11713 9199 11719 9225
rect 11745 9199 11751 9225
rect 13281 9199 13287 9225
rect 13313 9199 13319 9225
rect 13617 9199 13623 9225
rect 13649 9199 13655 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 10767 9193 10793 9199
rect 14911 9169 14937 9175
rect 11153 9143 11159 9169
rect 11185 9143 11191 9169
rect 11881 9143 11887 9169
rect 11913 9143 11919 9169
rect 14681 9143 14687 9169
rect 14713 9143 14719 9169
rect 14911 9137 14937 9143
rect 9535 9113 9561 9119
rect 6673 9087 6679 9113
rect 6705 9087 6711 9113
rect 9535 9081 9561 9087
rect 9983 9113 10009 9119
rect 9983 9081 10009 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 9871 8945 9897 8951
rect 7009 8919 7015 8945
rect 7041 8919 7047 8945
rect 9871 8913 9897 8919
rect 9927 8945 9953 8951
rect 11439 8945 11465 8951
rect 11265 8919 11271 8945
rect 11297 8919 11303 8945
rect 9927 8913 9953 8919
rect 11439 8913 11465 8919
rect 967 8889 993 8895
rect 10711 8889 10737 8895
rect 7625 8863 7631 8889
rect 7657 8863 7663 8889
rect 8689 8863 8695 8889
rect 8721 8863 8727 8889
rect 10929 8863 10935 8889
rect 10961 8863 10967 8889
rect 967 8857 993 8863
rect 10711 8857 10737 8863
rect 6735 8833 6761 8839
rect 9367 8833 9393 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 7065 8807 7071 8833
rect 7097 8807 7103 8833
rect 9025 8807 9031 8833
rect 9057 8807 9063 8833
rect 6735 8801 6761 8807
rect 9367 8801 9393 8807
rect 9647 8833 9673 8839
rect 10879 8833 10905 8839
rect 10201 8807 10207 8833
rect 10233 8807 10239 8833
rect 9647 8801 9673 8807
rect 10879 8801 10905 8807
rect 11551 8833 11577 8839
rect 11551 8801 11577 8807
rect 11719 8833 11745 8839
rect 11719 8801 11745 8807
rect 14071 8833 14097 8839
rect 14071 8801 14097 8807
rect 9591 8777 9617 8783
rect 6841 8751 6847 8777
rect 6873 8751 6879 8777
rect 9591 8745 9617 8751
rect 10039 8777 10065 8783
rect 10039 8745 10065 8751
rect 10319 8777 10345 8783
rect 10319 8745 10345 8751
rect 13903 8777 13929 8783
rect 13903 8745 13929 8751
rect 13959 8777 13985 8783
rect 13959 8745 13985 8751
rect 6791 8721 6817 8727
rect 6791 8689 6817 8695
rect 9535 8721 9561 8727
rect 9535 8689 9561 8695
rect 10263 8721 10289 8727
rect 11881 8695 11887 8721
rect 11913 8695 11919 8721
rect 10263 8689 10289 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 6623 8553 6649 8559
rect 11047 8553 11073 8559
rect 6953 8527 6959 8553
rect 6985 8527 6991 8553
rect 6623 8521 6649 8527
rect 11047 8521 11073 8527
rect 12615 8553 12641 8559
rect 12615 8521 12641 8527
rect 13231 8553 13257 8559
rect 13231 8521 13257 8527
rect 13343 8553 13369 8559
rect 13343 8521 13369 8527
rect 6847 8497 6873 8503
rect 11383 8497 11409 8503
rect 9081 8471 9087 8497
rect 9113 8471 9119 8497
rect 6847 8465 6873 8471
rect 11383 8465 11409 8471
rect 12951 8497 12977 8503
rect 12951 8465 12977 8471
rect 6567 8441 6593 8447
rect 2081 8415 2087 8441
rect 2113 8415 2119 8441
rect 6567 8409 6593 8415
rect 7015 8441 7041 8447
rect 10879 8441 10905 8447
rect 7121 8415 7127 8441
rect 7153 8415 7159 8441
rect 7849 8415 7855 8441
rect 7881 8415 7887 8441
rect 8745 8415 8751 8441
rect 8777 8415 8783 8441
rect 7015 8409 7041 8415
rect 10879 8409 10905 8415
rect 12671 8441 12697 8447
rect 12671 8409 12697 8415
rect 12783 8441 12809 8447
rect 12783 8409 12809 8415
rect 13567 8441 13593 8447
rect 13567 8409 13593 8415
rect 13735 8441 13761 8447
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 13735 8409 13761 8415
rect 7687 8385 7713 8391
rect 7687 8353 7713 8359
rect 7743 8385 7769 8391
rect 13287 8385 13313 8391
rect 10145 8359 10151 8385
rect 10177 8359 10183 8385
rect 19945 8359 19951 8385
rect 19977 8359 19983 8385
rect 7743 8353 7769 8359
rect 13287 8353 13313 8359
rect 967 8329 993 8335
rect 11439 8329 11465 8335
rect 7121 8303 7127 8329
rect 7153 8303 7159 8329
rect 967 8297 993 8303
rect 11439 8297 11465 8303
rect 13063 8329 13089 8335
rect 13063 8297 13089 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 7183 8161 7209 8167
rect 7183 8129 7209 8135
rect 14127 8161 14153 8167
rect 14127 8129 14153 8135
rect 7239 8105 7265 8111
rect 20007 8105 20033 8111
rect 1017 8079 1023 8105
rect 1049 8079 1055 8105
rect 4993 8079 4999 8105
rect 5025 8079 5031 8105
rect 6057 8079 6063 8105
rect 6089 8079 6095 8105
rect 12553 8079 12559 8105
rect 12585 8079 12591 8105
rect 13617 8079 13623 8105
rect 13649 8079 13655 8105
rect 7239 8073 7265 8079
rect 20007 8073 20033 8079
rect 8415 8049 8441 8055
rect 2137 8023 2143 8049
rect 2169 8023 2175 8049
rect 6393 8023 6399 8049
rect 6425 8023 6431 8049
rect 6841 8023 6847 8049
rect 6873 8023 6879 8049
rect 8415 8017 8441 8023
rect 8751 8049 8777 8055
rect 8751 8017 8777 8023
rect 10151 8049 10177 8055
rect 10151 8017 10177 8023
rect 11663 8049 11689 8055
rect 11663 8017 11689 8023
rect 11999 8049 12025 8055
rect 13735 8049 13761 8055
rect 12217 8023 12223 8049
rect 12249 8023 12255 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 11999 8017 12025 8023
rect 13735 8017 13761 8023
rect 8527 7993 8553 7999
rect 6729 7967 6735 7993
rect 6761 7967 6767 7993
rect 8527 7961 8553 7967
rect 10095 7993 10121 7999
rect 13847 7993 13873 7999
rect 11489 7967 11495 7993
rect 11521 7967 11527 7993
rect 11825 7967 11831 7993
rect 11857 7967 11863 7993
rect 10095 7961 10121 7967
rect 13847 7961 13873 7967
rect 13903 7993 13929 7999
rect 13903 7961 13929 7967
rect 14071 7993 14097 7999
rect 14071 7961 14097 7967
rect 8471 7937 8497 7943
rect 8471 7905 8497 7911
rect 9983 7937 10009 7943
rect 9983 7905 10009 7911
rect 14127 7937 14153 7943
rect 14127 7905 14153 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8751 7769 8777 7775
rect 8751 7737 8777 7743
rect 14407 7769 14433 7775
rect 14407 7737 14433 7743
rect 8863 7713 8889 7719
rect 7121 7687 7127 7713
rect 7153 7687 7159 7713
rect 8863 7681 8889 7687
rect 8919 7713 8945 7719
rect 9473 7687 9479 7713
rect 9505 7687 9511 7713
rect 11097 7687 11103 7713
rect 11129 7687 11135 7713
rect 13113 7687 13119 7713
rect 13145 7687 13151 7713
rect 8919 7681 8945 7687
rect 7457 7631 7463 7657
rect 7489 7631 7495 7657
rect 9081 7631 9087 7657
rect 9113 7631 9119 7657
rect 10761 7631 10767 7657
rect 10793 7631 10799 7657
rect 12721 7631 12727 7657
rect 12753 7631 12759 7657
rect 6057 7575 6063 7601
rect 6089 7575 6095 7601
rect 10537 7575 10543 7601
rect 10569 7575 10575 7601
rect 12161 7575 12167 7601
rect 12193 7575 12199 7601
rect 14177 7575 14183 7601
rect 14209 7575 14215 7601
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 12335 7321 12361 7327
rect 8185 7295 8191 7321
rect 8217 7295 8223 7321
rect 9249 7295 9255 7321
rect 9281 7295 9287 7321
rect 12335 7289 12361 7295
rect 7849 7239 7855 7265
rect 7881 7239 7887 7265
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 10929 1807 10935 1833
rect 10961 1807 10967 1833
rect 9311 1801 9337 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10369 1751 10375 1777
rect 10401 1751 10407 1777
rect 7855 1665 7881 1671
rect 7855 1633 7881 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9031 19111 9057 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 8527 18999 8553 19025
rect 10879 18999 10905 19025
rect 12279 18999 12305 19025
rect 9983 18943 10009 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 10039 18719 10065 18745
rect 13735 18719 13761 18745
rect 9535 18607 9561 18633
rect 13399 18607 13425 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 20119 18103 20145 18129
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 11663 14015 11689 14041
rect 11551 13903 11577 13929
rect 11719 13903 11745 13929
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9535 13567 9561 13593
rect 12111 13567 12137 13593
rect 8079 13511 8105 13537
rect 9815 13511 9841 13537
rect 10711 13511 10737 13537
rect 8471 13455 8497 13481
rect 9647 13455 9673 13481
rect 9759 13455 9785 13481
rect 11047 13455 11073 13481
rect 12335 13399 12361 13425
rect 20119 13399 20145 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8695 13231 8721 13257
rect 8807 13231 8833 13257
rect 11551 13231 11577 13257
rect 11831 13175 11857 13201
rect 8863 13119 8889 13145
rect 11271 13119 11297 13145
rect 11495 13119 11521 13145
rect 9871 13063 9897 13089
rect 10935 13063 10961 13089
rect 12671 13063 12697 13089
rect 11551 13007 11577 13033
rect 12615 13007 12641 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 10935 12839 10961 12865
rect 8359 12783 8385 12809
rect 12335 12783 12361 12809
rect 13399 12783 13425 12809
rect 6959 12727 6985 12753
rect 11943 12727 11969 12753
rect 7295 12671 7321 12697
rect 8583 12671 8609 12697
rect 8639 12671 8665 12697
rect 9031 12671 9057 12697
rect 9199 12671 9225 12697
rect 10655 12671 10681 12697
rect 10879 12671 10905 12697
rect 10991 12671 11017 12697
rect 11103 12671 11129 12697
rect 11159 12671 11185 12697
rect 8471 12615 8497 12641
rect 10767 12615 10793 12641
rect 13623 12615 13649 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8135 12447 8161 12473
rect 12167 12447 12193 12473
rect 12223 12447 12249 12473
rect 12279 12447 12305 12473
rect 2143 12335 2169 12361
rect 7071 12335 7097 12361
rect 7967 12335 7993 12361
rect 8135 12335 8161 12361
rect 8303 12335 8329 12361
rect 9031 12335 9057 12361
rect 11999 12335 12025 12361
rect 12111 12335 12137 12361
rect 5671 12279 5697 12305
rect 6735 12279 6761 12305
rect 9367 12279 9393 12305
rect 10431 12279 10457 12305
rect 967 12223 993 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 7519 11999 7545 12025
rect 9647 11999 9673 12025
rect 12727 11999 12753 12025
rect 12951 11999 12977 12025
rect 20007 11999 20033 12025
rect 7071 11943 7097 11969
rect 7463 11943 7489 11969
rect 7631 11943 7657 11969
rect 11271 11943 11297 11969
rect 18943 11943 18969 11969
rect 11663 11887 11689 11913
rect 13567 11887 13593 11913
rect 7015 11831 7041 11857
rect 7127 11831 7153 11857
rect 7239 11831 7265 11857
rect 9479 11831 9505 11857
rect 9591 11831 9617 11857
rect 9703 11831 9729 11857
rect 13623 11831 13649 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 10879 11663 10905 11689
rect 11159 11663 11185 11689
rect 11719 11663 11745 11689
rect 12727 11663 12753 11689
rect 8807 11607 8833 11633
rect 8919 11607 8945 11633
rect 9199 11607 9225 11633
rect 10487 11607 10513 11633
rect 12671 11607 12697 11633
rect 12951 11607 12977 11633
rect 13679 11607 13705 11633
rect 6959 11551 6985 11577
rect 9255 11551 9281 11577
rect 9927 11551 9953 11577
rect 10319 11551 10345 11577
rect 10599 11551 10625 11577
rect 10767 11551 10793 11577
rect 11047 11551 11073 11577
rect 12783 11551 12809 11577
rect 13343 11551 13369 11577
rect 18831 11551 18857 11577
rect 7351 11495 7377 11521
rect 8415 11495 8441 11521
rect 8863 11495 8889 11521
rect 10823 11495 10849 11521
rect 11663 11495 11689 11521
rect 14743 11495 14769 11521
rect 14967 11495 14993 11521
rect 9199 11439 9225 11465
rect 9871 11439 9897 11465
rect 11215 11439 11241 11465
rect 11831 11439 11857 11465
rect 13063 11439 13089 11465
rect 13119 11439 13145 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 967 11215 993 11241
rect 8191 11215 8217 11241
rect 11887 11215 11913 11241
rect 20007 11215 20033 11241
rect 2143 11159 2169 11185
rect 6847 11159 6873 11185
rect 6959 11159 6985 11185
rect 7183 11159 7209 11185
rect 8303 11159 8329 11185
rect 8359 11159 8385 11185
rect 10039 11159 10065 11185
rect 10263 11159 10289 11185
rect 11215 11159 11241 11185
rect 11495 11159 11521 11185
rect 11775 11159 11801 11185
rect 11999 11159 12025 11185
rect 12279 11159 12305 11185
rect 13175 11159 13201 11185
rect 13343 11159 13369 11185
rect 13623 11159 13649 11185
rect 13679 11159 13705 11185
rect 14239 11159 14265 11185
rect 18831 11159 18857 11185
rect 8135 11103 8161 11129
rect 9143 11103 9169 11129
rect 9311 11103 9337 11129
rect 9759 11103 9785 11129
rect 9871 11103 9897 11129
rect 10375 11103 10401 11129
rect 11663 11103 11689 11129
rect 13455 11103 13481 11129
rect 14295 11103 14321 11129
rect 6903 11047 6929 11073
rect 8807 11047 8833 11073
rect 8975 11047 9001 11073
rect 9535 11047 9561 11073
rect 10711 11047 10737 11073
rect 10879 11047 10905 11073
rect 11103 11047 11129 11073
rect 11775 11047 11801 11073
rect 12167 11047 12193 11073
rect 13287 11047 13313 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8807 10879 8833 10905
rect 9311 10879 9337 10905
rect 8359 10823 8385 10849
rect 8975 10823 9001 10849
rect 6903 10767 6929 10793
rect 7071 10767 7097 10793
rect 7239 10767 7265 10793
rect 7407 10767 7433 10793
rect 9199 10767 9225 10793
rect 9535 10767 9561 10793
rect 9759 10767 9785 10793
rect 12615 10767 12641 10793
rect 5447 10711 5473 10737
rect 6511 10711 6537 10737
rect 7295 10711 7321 10737
rect 11719 10711 11745 10737
rect 15023 10711 15049 10737
rect 8415 10655 8441 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 6735 10487 6761 10513
rect 6903 10487 6929 10513
rect 967 10431 993 10457
rect 4999 10431 5025 10457
rect 9031 10431 9057 10457
rect 11775 10431 11801 10457
rect 12615 10431 12641 10457
rect 20007 10431 20033 10457
rect 2143 10375 2169 10401
rect 6455 10375 6481 10401
rect 10039 10375 10065 10401
rect 10767 10375 10793 10401
rect 10935 10375 10961 10401
rect 11383 10375 11409 10401
rect 11887 10375 11913 10401
rect 12391 10375 12417 10401
rect 12839 10375 12865 10401
rect 18831 10375 18857 10401
rect 6063 10319 6089 10345
rect 6791 10319 6817 10345
rect 11159 10319 11185 10345
rect 11439 10319 11465 10345
rect 12167 10319 12193 10345
rect 12503 10319 12529 10345
rect 12671 10319 12697 10345
rect 13007 10319 13033 10345
rect 13511 10319 13537 10345
rect 13567 10319 13593 10345
rect 10711 10263 10737 10289
rect 13679 10263 13705 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 10263 10095 10289 10121
rect 10991 10095 11017 10121
rect 11103 10095 11129 10121
rect 11943 10095 11969 10121
rect 6567 10039 6593 10065
rect 6679 10039 6705 10065
rect 6847 10039 6873 10065
rect 6903 10039 6929 10065
rect 9087 10039 9113 10065
rect 10375 10039 10401 10065
rect 11159 10039 11185 10065
rect 11887 10039 11913 10065
rect 11999 10039 12025 10065
rect 12671 10039 12697 10065
rect 12727 10067 12753 10093
rect 12895 10039 12921 10065
rect 13735 10039 13761 10065
rect 2143 9983 2169 10009
rect 6511 9983 6537 10009
rect 9423 9983 9449 10009
rect 9591 9983 9617 10009
rect 10319 9983 10345 10009
rect 13007 9983 13033 10009
rect 13231 9983 13257 10009
rect 13343 9983 13369 10009
rect 9143 9927 9169 9953
rect 9871 9927 9897 9953
rect 13119 9927 13145 9953
rect 14799 9927 14825 9953
rect 15023 9927 15049 9953
rect 967 9871 993 9897
rect 6847 9871 6873 9897
rect 8975 9871 9001 9897
rect 9535 9871 9561 9897
rect 12671 9871 12697 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 11215 9703 11241 9729
rect 11943 9703 11969 9729
rect 967 9647 993 9673
rect 4999 9647 5025 9673
rect 9367 9647 9393 9673
rect 13231 9647 13257 9673
rect 14295 9647 14321 9673
rect 2143 9591 2169 9617
rect 6455 9591 6481 9617
rect 8807 9591 8833 9617
rect 9423 9591 9449 9617
rect 9591 9591 9617 9617
rect 10039 9591 10065 9617
rect 11663 9591 11689 9617
rect 12895 9591 12921 9617
rect 14575 9591 14601 9617
rect 14687 9591 14713 9617
rect 6063 9535 6089 9561
rect 6903 9535 6929 9561
rect 7071 9535 7097 9561
rect 9199 9535 9225 9561
rect 11271 9535 11297 9561
rect 8975 9479 9001 9505
rect 9871 9479 9897 9505
rect 11775 9479 11801 9505
rect 11887 9479 11913 9505
rect 14631 9479 14657 9505
rect 14799 9479 14825 9505
rect 15079 9479 15105 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 5895 9311 5921 9337
rect 6511 9311 6537 9337
rect 9815 9311 9841 9337
rect 6399 9255 6425 9281
rect 7127 9255 7153 9281
rect 9759 9255 9785 9281
rect 10151 9255 10177 9281
rect 10879 9255 10905 9281
rect 10935 9255 10961 9281
rect 11551 9255 11577 9281
rect 5839 9199 5865 9225
rect 6567 9199 6593 9225
rect 6791 9199 6817 9225
rect 7295 9199 7321 9225
rect 9255 9199 9281 9225
rect 9423 9199 9449 9225
rect 9647 9199 9673 9225
rect 10039 9199 10065 9225
rect 10319 9199 10345 9225
rect 10375 9199 10401 9225
rect 10431 9199 10457 9225
rect 10767 9199 10793 9225
rect 11327 9199 11353 9225
rect 11719 9199 11745 9225
rect 13287 9199 13313 9225
rect 13623 9199 13649 9225
rect 18831 9199 18857 9225
rect 11159 9143 11185 9169
rect 11887 9143 11913 9169
rect 14687 9143 14713 9169
rect 14911 9143 14937 9169
rect 6679 9087 6705 9113
rect 9535 9087 9561 9113
rect 9983 9087 10009 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 7015 8919 7041 8945
rect 9871 8919 9897 8945
rect 9927 8919 9953 8945
rect 11271 8919 11297 8945
rect 11439 8919 11465 8945
rect 967 8863 993 8889
rect 7631 8863 7657 8889
rect 8695 8863 8721 8889
rect 10711 8863 10737 8889
rect 10935 8863 10961 8889
rect 2143 8807 2169 8833
rect 6735 8807 6761 8833
rect 7071 8807 7097 8833
rect 9031 8807 9057 8833
rect 9367 8807 9393 8833
rect 9647 8807 9673 8833
rect 10207 8807 10233 8833
rect 10879 8807 10905 8833
rect 11551 8807 11577 8833
rect 11719 8807 11745 8833
rect 14071 8807 14097 8833
rect 6847 8751 6873 8777
rect 9591 8751 9617 8777
rect 10039 8751 10065 8777
rect 10319 8751 10345 8777
rect 13903 8751 13929 8777
rect 13959 8751 13985 8777
rect 6791 8695 6817 8721
rect 9535 8695 9561 8721
rect 10263 8695 10289 8721
rect 11887 8695 11913 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 6623 8527 6649 8553
rect 6959 8527 6985 8553
rect 11047 8527 11073 8553
rect 12615 8527 12641 8553
rect 13231 8527 13257 8553
rect 13343 8527 13369 8553
rect 6847 8471 6873 8497
rect 9087 8471 9113 8497
rect 11383 8471 11409 8497
rect 12951 8471 12977 8497
rect 2087 8415 2113 8441
rect 6567 8415 6593 8441
rect 7015 8415 7041 8441
rect 7127 8415 7153 8441
rect 7855 8415 7881 8441
rect 8751 8415 8777 8441
rect 10879 8415 10905 8441
rect 12671 8415 12697 8441
rect 12783 8415 12809 8441
rect 13567 8415 13593 8441
rect 13735 8415 13761 8441
rect 18831 8415 18857 8441
rect 7687 8359 7713 8385
rect 7743 8359 7769 8385
rect 10151 8359 10177 8385
rect 13287 8359 13313 8385
rect 19951 8359 19977 8385
rect 967 8303 993 8329
rect 7127 8303 7153 8329
rect 11439 8303 11465 8329
rect 13063 8303 13089 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 7183 8135 7209 8161
rect 14127 8135 14153 8161
rect 1023 8079 1049 8105
rect 4999 8079 5025 8105
rect 6063 8079 6089 8105
rect 7239 8079 7265 8105
rect 12559 8079 12585 8105
rect 13623 8079 13649 8105
rect 20007 8079 20033 8105
rect 2143 8023 2169 8049
rect 6399 8023 6425 8049
rect 6847 8023 6873 8049
rect 8415 8023 8441 8049
rect 8751 8023 8777 8049
rect 10151 8023 10177 8049
rect 11663 8023 11689 8049
rect 11999 8023 12025 8049
rect 12223 8023 12249 8049
rect 13735 8023 13761 8049
rect 18831 8023 18857 8049
rect 6735 7967 6761 7993
rect 8527 7967 8553 7993
rect 10095 7967 10121 7993
rect 11495 7967 11521 7993
rect 11831 7967 11857 7993
rect 13847 7967 13873 7993
rect 13903 7967 13929 7993
rect 14071 7967 14097 7993
rect 8471 7911 8497 7937
rect 9983 7911 10009 7937
rect 14127 7911 14153 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8751 7743 8777 7769
rect 14407 7743 14433 7769
rect 7127 7687 7153 7713
rect 8863 7687 8889 7713
rect 8919 7687 8945 7713
rect 9479 7687 9505 7713
rect 11103 7687 11129 7713
rect 13119 7687 13145 7713
rect 7463 7631 7489 7657
rect 9087 7631 9113 7657
rect 10767 7631 10793 7657
rect 12727 7631 12753 7657
rect 6063 7575 6089 7601
rect 10543 7575 10569 7601
rect 12167 7575 12193 7601
rect 14183 7575 14209 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 8191 7295 8217 7321
rect 9255 7295 9281 7321
rect 12335 7295 12361 7321
rect 7855 7239 7881 7265
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 10935 1807 10961 1833
rect 8807 1751 8833 1777
rect 10375 1751 10401 1777
rect 7855 1639 7881 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 9408 20600 9464 21000
rect 9744 20600 9800 21000
rect 11088 20600 11144 21000
rect 11760 20600 11816 21000
rect 13104 20600 13160 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8414 19138 8442 20600
rect 8414 19105 8442 19110
rect 9030 19138 9058 19143
rect 9030 19091 9058 19110
rect 8526 19025 8554 19031
rect 8526 18999 8527 19025
rect 8553 18999 8554 19025
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8526 15974 8554 18999
rect 9422 18746 9450 20600
rect 9758 19810 9786 20600
rect 9758 19782 10010 19810
rect 9982 18969 10010 19782
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 11774 19138 11802 20600
rect 11774 19105 11802 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 9982 18943 9983 18969
rect 10009 18943 10010 18969
rect 9982 18937 10010 18943
rect 10878 19025 10906 19031
rect 10878 18999 10879 19025
rect 10905 18999 10906 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9422 18713 9450 18718
rect 10038 18746 10066 18751
rect 10038 18699 10066 18718
rect 8414 15946 8554 15974
rect 9534 18633 9562 18639
rect 9534 18607 9535 18633
rect 9561 18607 9562 18633
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 6958 13538 6986 13543
rect 2086 13482 2114 13487
rect 966 12250 994 12255
rect 966 12203 994 12222
rect 966 11242 994 11247
rect 966 11195 994 11214
rect 2086 10794 2114 13454
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 6958 12754 6986 13510
rect 8078 13538 8106 13543
rect 8078 13491 8106 13510
rect 8414 13454 8442 15946
rect 9534 13594 9562 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9534 13593 9786 13594
rect 9534 13567 9535 13593
rect 9561 13567 9786 13593
rect 9534 13566 9786 13567
rect 9534 13561 9562 13566
rect 9198 13538 9226 13543
rect 8358 13426 8442 13454
rect 8470 13481 8498 13487
rect 8470 13455 8471 13481
rect 8497 13455 8498 13481
rect 8470 13454 8498 13455
rect 8806 13482 8834 13487
rect 8470 13426 8722 13454
rect 8358 12810 8386 13426
rect 8694 13257 8722 13426
rect 8694 13231 8695 13257
rect 8721 13231 8722 13257
rect 8694 13225 8722 13231
rect 8806 13257 8834 13454
rect 8806 13231 8807 13257
rect 8833 13231 8834 13257
rect 8806 13225 8834 13231
rect 8862 13146 8890 13151
rect 8862 13145 9114 13146
rect 8862 13119 8863 13145
rect 8889 13119 9114 13145
rect 8862 13118 9114 13119
rect 8862 13113 8890 13118
rect 8358 12809 8610 12810
rect 8358 12783 8359 12809
rect 8385 12783 8610 12809
rect 8358 12782 8610 12783
rect 8358 12777 8386 12782
rect 6958 12753 7098 12754
rect 6958 12727 6959 12753
rect 6985 12727 7098 12753
rect 6958 12726 7098 12727
rect 6958 12721 6986 12726
rect 2142 12362 2170 12367
rect 2142 12315 2170 12334
rect 5670 12362 5698 12367
rect 7070 12362 7098 12726
rect 7294 12697 7322 12703
rect 7294 12671 7295 12697
rect 7321 12671 7322 12697
rect 7294 12474 7322 12671
rect 8582 12697 8610 12782
rect 9086 12754 9114 13118
rect 9086 12726 9170 12754
rect 8582 12671 8583 12697
rect 8609 12671 8610 12697
rect 8582 12665 8610 12671
rect 8638 12698 8666 12703
rect 9030 12698 9058 12703
rect 8638 12697 9114 12698
rect 8638 12671 8639 12697
rect 8665 12671 9031 12697
rect 9057 12671 9114 12697
rect 8638 12670 9114 12671
rect 8638 12665 8666 12670
rect 9030 12665 9058 12670
rect 8470 12642 8498 12647
rect 8302 12641 8498 12642
rect 8302 12615 8471 12641
rect 8497 12615 8498 12641
rect 8302 12614 8498 12615
rect 7294 12441 7322 12446
rect 8134 12474 8162 12479
rect 8134 12427 8162 12446
rect 7966 12362 7994 12367
rect 5670 12305 5698 12334
rect 6958 12361 7098 12362
rect 6958 12335 7071 12361
rect 7097 12335 7098 12361
rect 6958 12334 7098 12335
rect 5670 12279 5671 12305
rect 5697 12279 5698 12305
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 5670 11858 5698 12279
rect 6734 12306 6762 12311
rect 6734 12259 6762 12278
rect 5670 11825 5698 11830
rect 6958 11578 6986 12334
rect 7070 12329 7098 12334
rect 7630 12361 7994 12362
rect 7630 12335 7967 12361
rect 7993 12335 7994 12361
rect 7630 12334 7994 12335
rect 7518 12306 7546 12311
rect 7518 12025 7546 12278
rect 7518 11999 7519 12025
rect 7545 11999 7546 12025
rect 7518 11993 7546 11999
rect 7070 11970 7098 11975
rect 7462 11970 7490 11975
rect 7070 11969 7490 11970
rect 7070 11943 7071 11969
rect 7097 11943 7463 11969
rect 7489 11943 7490 11969
rect 7070 11942 7490 11943
rect 7070 11937 7098 11942
rect 7462 11937 7490 11942
rect 7630 11969 7658 12334
rect 7966 12329 7994 12334
rect 8134 12361 8162 12367
rect 8134 12335 8135 12361
rect 8161 12335 8162 12361
rect 7630 11943 7631 11969
rect 7657 11943 7658 11969
rect 7014 11858 7042 11863
rect 7126 11858 7154 11863
rect 7014 11857 7098 11858
rect 7014 11831 7015 11857
rect 7041 11831 7098 11857
rect 7014 11830 7098 11831
rect 7014 11825 7042 11830
rect 6958 11577 7042 11578
rect 6958 11551 6959 11577
rect 6985 11551 7042 11577
rect 6958 11550 7042 11551
rect 6958 11545 6986 11550
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 6846 11298 6874 11303
rect 2142 11186 2170 11191
rect 2142 11139 2170 11158
rect 5446 11186 5474 11191
rect 2086 10761 2114 10766
rect 5446 10737 5474 11158
rect 6846 11185 6874 11270
rect 6846 11159 6847 11185
rect 6873 11159 6874 11185
rect 6846 11153 6874 11159
rect 6958 11186 6986 11191
rect 6958 11139 6986 11158
rect 6902 11073 6930 11079
rect 6902 11047 6903 11073
rect 6929 11047 6930 11073
rect 6902 10906 6930 11047
rect 6846 10878 6930 10906
rect 5446 10711 5447 10737
rect 5473 10711 5474 10737
rect 5446 10705 5474 10711
rect 6454 10738 6482 10743
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 966 10457 994 10463
rect 966 10431 967 10457
rect 993 10431 994 10457
rect 966 10122 994 10431
rect 4998 10458 5026 10463
rect 4998 10411 5026 10430
rect 2142 10402 2170 10407
rect 2142 10355 2170 10374
rect 6454 10401 6482 10710
rect 6510 10738 6538 10743
rect 6510 10737 6762 10738
rect 6510 10711 6511 10737
rect 6537 10711 6762 10737
rect 6510 10710 6762 10711
rect 6510 10705 6538 10710
rect 6734 10513 6762 10710
rect 6734 10487 6735 10513
rect 6761 10487 6762 10513
rect 6734 10481 6762 10487
rect 6846 10514 6874 10878
rect 6902 10794 6930 10799
rect 7014 10794 7042 11550
rect 7070 11298 7098 11830
rect 7126 11811 7154 11830
rect 7238 11857 7266 11863
rect 7238 11831 7239 11857
rect 7265 11831 7266 11857
rect 7238 11634 7266 11831
rect 7070 11265 7098 11270
rect 7182 11606 7238 11634
rect 7182 11185 7210 11606
rect 7238 11601 7266 11606
rect 7350 11522 7378 11527
rect 7350 11475 7378 11494
rect 7182 11159 7183 11185
rect 7209 11159 7210 11185
rect 7182 11153 7210 11159
rect 7630 11186 7658 11943
rect 7630 11153 7658 11158
rect 8134 11130 8162 12335
rect 8302 12361 8330 12614
rect 8470 12609 8498 12614
rect 8302 12335 8303 12361
rect 8329 12335 8330 12361
rect 8302 12329 8330 12335
rect 9030 12361 9058 12367
rect 9030 12335 9031 12361
rect 9057 12335 9058 12361
rect 8302 11690 8330 11695
rect 8190 11522 8218 11527
rect 8190 11241 8218 11494
rect 8190 11215 8191 11241
rect 8217 11215 8218 11241
rect 8190 11209 8218 11215
rect 8302 11185 8330 11662
rect 8806 11690 8834 11695
rect 8806 11633 8834 11662
rect 8806 11607 8807 11633
rect 8833 11607 8834 11633
rect 8806 11601 8834 11607
rect 8918 11633 8946 11639
rect 8918 11607 8919 11633
rect 8945 11607 8946 11633
rect 8414 11522 8442 11527
rect 8414 11521 8498 11522
rect 8414 11495 8415 11521
rect 8441 11495 8498 11521
rect 8414 11494 8498 11495
rect 8414 11489 8442 11494
rect 8302 11159 8303 11185
rect 8329 11159 8330 11185
rect 8302 11153 8330 11159
rect 8358 11186 8386 11191
rect 8358 11139 8386 11158
rect 8134 11083 8162 11102
rect 7238 11018 7266 11023
rect 6902 10793 7042 10794
rect 6902 10767 6903 10793
rect 6929 10767 7042 10793
rect 6902 10766 7042 10767
rect 7070 10793 7098 10799
rect 7070 10767 7071 10793
rect 7097 10767 7098 10793
rect 6902 10738 6930 10766
rect 6902 10705 6930 10710
rect 6902 10514 6930 10519
rect 6846 10513 6930 10514
rect 6846 10487 6903 10513
rect 6929 10487 6930 10513
rect 6846 10486 6930 10487
rect 6902 10481 6930 10486
rect 6454 10375 6455 10401
rect 6481 10375 6482 10401
rect 966 10089 994 10094
rect 6062 10345 6090 10351
rect 6062 10319 6063 10345
rect 6089 10319 6090 10345
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 6062 9898 6090 10319
rect 6454 10094 6482 10375
rect 6062 9865 6090 9870
rect 6398 10066 6482 10094
rect 6566 10458 6594 10463
rect 7070 10458 7098 10767
rect 7238 10793 7266 10990
rect 8470 10906 8498 11494
rect 8862 11521 8890 11527
rect 8862 11495 8863 11521
rect 8889 11495 8890 11521
rect 8358 10878 8470 10906
rect 8358 10849 8386 10878
rect 8470 10859 8498 10878
rect 8526 11466 8554 11471
rect 8526 11130 8554 11438
rect 8862 11186 8890 11495
rect 8862 11153 8890 11158
rect 8358 10823 8359 10849
rect 8385 10823 8386 10849
rect 8358 10817 8386 10823
rect 7238 10767 7239 10793
rect 7265 10767 7266 10793
rect 7238 10761 7266 10767
rect 7406 10793 7434 10799
rect 8526 10794 8554 11102
rect 8918 11130 8946 11607
rect 8918 11097 8946 11102
rect 8974 11578 9002 11583
rect 8806 11074 8834 11079
rect 8974 11074 9002 11550
rect 8806 11073 8890 11074
rect 8806 11047 8807 11073
rect 8833 11047 8890 11073
rect 8806 11046 8890 11047
rect 8806 11041 8834 11046
rect 8806 10906 8834 10911
rect 8806 10859 8834 10878
rect 7406 10767 7407 10793
rect 7433 10767 7434 10793
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 966 9673 994 9679
rect 966 9647 967 9673
rect 993 9647 994 9673
rect 966 9450 994 9647
rect 4998 9674 5026 9679
rect 6398 9674 6426 10066
rect 6566 10065 6594 10430
rect 6958 10430 7098 10458
rect 7294 10737 7322 10743
rect 7294 10711 7295 10737
rect 7321 10711 7322 10737
rect 6958 10402 6986 10430
rect 6790 10374 6986 10402
rect 6790 10345 6818 10374
rect 6790 10319 6791 10345
rect 6817 10319 6818 10345
rect 6566 10039 6567 10065
rect 6593 10039 6594 10065
rect 6566 10033 6594 10039
rect 6678 10066 6706 10071
rect 6678 10019 6706 10038
rect 6510 10009 6538 10015
rect 6510 9983 6511 10009
rect 6537 9983 6538 10009
rect 4998 9627 5026 9646
rect 6342 9646 6482 9674
rect 2142 9618 2170 9623
rect 2142 9571 2170 9590
rect 6062 9562 6090 9567
rect 966 9417 994 9422
rect 5894 9561 6090 9562
rect 5894 9535 6063 9561
rect 6089 9535 6090 9561
rect 5894 9534 6090 9535
rect 5838 9338 5866 9343
rect 5838 9225 5866 9310
rect 5894 9337 5922 9534
rect 6062 9529 6090 9534
rect 5894 9311 5895 9337
rect 5921 9311 5922 9337
rect 5894 9305 5922 9311
rect 5838 9199 5839 9225
rect 5865 9199 5866 9225
rect 5838 9193 5866 9199
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8889 994 8895
rect 966 8863 967 8889
rect 993 8863 994 8889
rect 966 8442 994 8863
rect 2142 8833 2170 8839
rect 2142 8807 2143 8833
rect 2169 8807 2170 8833
rect 966 8409 994 8414
rect 2086 8441 2114 8447
rect 2086 8415 2087 8441
rect 2113 8415 2114 8441
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 966 8073 994 8078
rect 1022 8105 1050 8111
rect 1022 8079 1023 8105
rect 1049 8079 1050 8105
rect 1022 7770 1050 8079
rect 2086 7994 2114 8415
rect 2142 8330 2170 8807
rect 6062 8722 6090 8727
rect 2142 8297 2170 8302
rect 4998 8330 5026 8335
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 4998 8105 5026 8302
rect 4998 8079 4999 8105
rect 5025 8079 5026 8105
rect 4998 8073 5026 8079
rect 6062 8105 6090 8694
rect 6062 8079 6063 8105
rect 6089 8079 6090 8105
rect 6062 8073 6090 8079
rect 2142 8050 2170 8055
rect 2142 8003 2170 8022
rect 6006 8050 6034 8055
rect 6342 8050 6370 9646
rect 6454 9617 6482 9646
rect 6454 9591 6455 9617
rect 6481 9591 6482 9617
rect 6454 9585 6482 9591
rect 6510 9506 6538 9983
rect 6398 9478 6538 9506
rect 6566 9674 6594 9679
rect 6790 9674 6818 10319
rect 7294 10094 7322 10711
rect 6846 10066 6874 10071
rect 6846 10019 6874 10038
rect 6902 10066 7322 10094
rect 7406 10290 7434 10767
rect 8470 10766 8554 10794
rect 6902 10065 6930 10066
rect 6902 10039 6903 10065
rect 6929 10039 6930 10065
rect 6902 10033 6930 10039
rect 6846 9898 6874 9903
rect 6846 9851 6874 9870
rect 6790 9646 7098 9674
rect 6398 9281 6426 9478
rect 6510 9338 6538 9357
rect 6510 9305 6538 9310
rect 6398 9255 6399 9281
rect 6425 9255 6426 9281
rect 6398 9226 6426 9255
rect 6398 9193 6426 9198
rect 6566 9225 6594 9646
rect 6902 9561 6930 9567
rect 6902 9535 6903 9561
rect 6929 9535 6930 9561
rect 6566 9199 6567 9225
rect 6593 9199 6594 9225
rect 6566 9193 6594 9199
rect 6734 9226 6762 9231
rect 6678 9113 6706 9119
rect 6678 9087 6679 9113
rect 6705 9087 6706 9113
rect 6678 8946 6706 9087
rect 6678 8913 6706 8918
rect 6734 8890 6762 9198
rect 6790 9226 6818 9231
rect 6902 9226 6930 9535
rect 6790 9225 6930 9226
rect 6790 9199 6791 9225
rect 6817 9199 6930 9225
rect 6790 9198 6930 9199
rect 6790 9193 6818 9198
rect 6902 9114 6930 9198
rect 6902 9081 6930 9086
rect 7070 9561 7098 9646
rect 7070 9535 7071 9561
rect 7097 9535 7098 9561
rect 7014 8946 7042 8951
rect 7014 8899 7042 8918
rect 6734 8862 6930 8890
rect 6734 8833 6762 8862
rect 6734 8807 6735 8833
rect 6761 8807 6762 8833
rect 6734 8801 6762 8807
rect 6846 8777 6874 8783
rect 6846 8751 6847 8777
rect 6873 8751 6874 8777
rect 6790 8722 6818 8727
rect 6790 8675 6818 8694
rect 6846 8610 6874 8751
rect 6622 8582 6874 8610
rect 6622 8553 6650 8582
rect 6622 8527 6623 8553
rect 6649 8527 6650 8553
rect 6622 8521 6650 8527
rect 6846 8498 6874 8503
rect 6902 8498 6930 8862
rect 7070 8834 7098 9535
rect 7126 9281 7154 9287
rect 7126 9255 7127 9281
rect 7153 9255 7154 9281
rect 7126 9226 7154 9255
rect 7126 9193 7154 9198
rect 7294 9225 7322 9231
rect 7294 9199 7295 9225
rect 7321 9199 7322 9225
rect 7070 8833 7154 8834
rect 7070 8807 7071 8833
rect 7097 8807 7154 8833
rect 7070 8806 7154 8807
rect 7070 8801 7098 8806
rect 6846 8497 6930 8498
rect 6846 8471 6847 8497
rect 6873 8471 6930 8497
rect 6846 8470 6930 8471
rect 6958 8553 6986 8559
rect 6958 8527 6959 8553
rect 6985 8527 6986 8553
rect 6846 8465 6874 8470
rect 6566 8441 6594 8447
rect 6566 8415 6567 8441
rect 6593 8415 6594 8441
rect 6566 8330 6594 8415
rect 6566 8297 6594 8302
rect 6846 8330 6874 8335
rect 6398 8050 6426 8055
rect 6342 8022 6398 8050
rect 2086 7961 2114 7966
rect 1022 7737 1050 7742
rect 6006 7602 6034 8022
rect 6398 8003 6426 8022
rect 6846 8049 6874 8302
rect 6846 8023 6847 8049
rect 6873 8023 6874 8049
rect 6846 8017 6874 8023
rect 6958 8050 6986 8527
rect 7014 8441 7042 8447
rect 7014 8415 7015 8441
rect 7041 8415 7042 8441
rect 7014 8218 7042 8415
rect 7126 8441 7154 8806
rect 7294 8498 7322 9199
rect 7406 8946 7434 10262
rect 8414 10681 8442 10687
rect 8414 10655 8415 10681
rect 8441 10655 8442 10681
rect 7406 8913 7434 8918
rect 7630 10010 7658 10015
rect 7630 9226 7658 9982
rect 8414 9898 8442 10655
rect 8414 9865 8442 9870
rect 7630 8889 7658 9198
rect 7630 8863 7631 8889
rect 7657 8863 7658 8889
rect 7630 8857 7658 8863
rect 7294 8465 7322 8470
rect 7686 8498 7714 8503
rect 7126 8415 7127 8441
rect 7153 8415 7154 8441
rect 7126 8409 7154 8415
rect 7686 8385 7714 8470
rect 7854 8441 7882 8447
rect 7854 8415 7855 8441
rect 7881 8415 7882 8441
rect 7686 8359 7687 8385
rect 7713 8359 7714 8385
rect 7686 8353 7714 8359
rect 7742 8386 7770 8391
rect 7742 8339 7770 8358
rect 7126 8330 7154 8335
rect 7126 8283 7154 8302
rect 7014 8190 7210 8218
rect 7182 8161 7210 8190
rect 7182 8135 7183 8161
rect 7209 8135 7210 8161
rect 7182 8129 7210 8135
rect 7238 8106 7266 8111
rect 7238 8059 7266 8078
rect 7462 8050 7490 8055
rect 6958 8022 7154 8050
rect 6734 7994 6762 7999
rect 6734 7947 6762 7966
rect 7126 7713 7154 8022
rect 7126 7687 7127 7713
rect 7153 7687 7154 7713
rect 7126 7681 7154 7687
rect 7462 7658 7490 8022
rect 7854 7994 7882 8415
rect 8414 8050 8442 8055
rect 8470 8050 8498 10766
rect 8806 9954 8834 9959
rect 8806 9617 8834 9926
rect 8862 9898 8890 11046
rect 8974 11027 9002 11046
rect 8974 10850 9002 10855
rect 8974 10803 9002 10822
rect 9030 10457 9058 12335
rect 9030 10431 9031 10457
rect 9057 10431 9058 10457
rect 8974 9898 9002 9903
rect 8862 9870 8974 9898
rect 8974 9851 9002 9870
rect 9030 9842 9058 10431
rect 9086 10402 9114 12670
rect 9142 11858 9170 12726
rect 9198 12697 9226 13510
rect 9646 13482 9674 13487
rect 9646 13435 9674 13454
rect 9758 13481 9786 13566
rect 9814 13538 9842 13543
rect 9814 13491 9842 13510
rect 10710 13537 10738 13543
rect 10710 13511 10711 13537
rect 10737 13511 10738 13537
rect 9758 13455 9759 13481
rect 9785 13455 9786 13481
rect 9758 13449 9786 13455
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10710 13202 10738 13511
rect 10710 13169 10738 13174
rect 10878 13202 10906 18999
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 12278 15974 12306 18999
rect 13118 18746 13146 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 13118 18713 13146 18718
rect 13734 18746 13762 18751
rect 13734 18699 13762 18718
rect 12110 15946 12306 15974
rect 13398 18633 13426 18639
rect 13398 18607 13399 18633
rect 13425 18607 13426 18633
rect 11662 14042 11690 14047
rect 11662 13995 11690 14014
rect 12110 14042 12138 15946
rect 11550 13929 11578 13935
rect 11550 13903 11551 13929
rect 11577 13903 11578 13929
rect 11046 13482 11074 13487
rect 11046 13481 11466 13482
rect 11046 13455 11047 13481
rect 11073 13455 11466 13481
rect 11046 13454 11466 13455
rect 11046 13449 11074 13454
rect 11158 13314 11186 13319
rect 10878 13174 11074 13202
rect 10822 13146 10850 13151
rect 9870 13090 9898 13095
rect 9870 13043 9898 13062
rect 9198 12671 9199 12697
rect 9225 12671 9226 12697
rect 9198 12665 9226 12671
rect 10654 12698 10682 12703
rect 10654 12651 10682 12670
rect 10822 12698 10850 13118
rect 10878 13090 10906 13174
rect 10878 13057 10906 13062
rect 10934 13089 10962 13095
rect 10934 13063 10935 13089
rect 10961 13063 10962 13089
rect 10934 12865 10962 13063
rect 10934 12839 10935 12865
rect 10961 12839 10962 12865
rect 10934 12833 10962 12839
rect 10878 12698 10906 12703
rect 10822 12697 10906 12698
rect 10822 12671 10879 12697
rect 10905 12671 10906 12697
rect 10822 12670 10906 12671
rect 10766 12642 10794 12647
rect 10710 12641 10794 12642
rect 10710 12615 10767 12641
rect 10793 12615 10794 12641
rect 10710 12614 10794 12615
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9366 12306 9394 12311
rect 10430 12306 10458 12311
rect 9366 12305 9674 12306
rect 9366 12279 9367 12305
rect 9393 12279 9674 12305
rect 9366 12278 9674 12279
rect 9366 12273 9394 12278
rect 9646 12025 9674 12278
rect 9646 11999 9647 12025
rect 9673 11999 9674 12025
rect 9646 11993 9674 11999
rect 10318 12305 10458 12306
rect 10318 12279 10431 12305
rect 10457 12279 10458 12305
rect 10318 12278 10458 12279
rect 9478 11858 9506 11863
rect 9142 11857 9562 11858
rect 9142 11831 9479 11857
rect 9505 11831 9562 11857
rect 9142 11830 9562 11831
rect 9478 11825 9506 11830
rect 9198 11634 9226 11639
rect 9142 11633 9226 11634
rect 9142 11607 9199 11633
rect 9225 11607 9226 11633
rect 9142 11606 9226 11607
rect 9142 11354 9170 11606
rect 9198 11601 9226 11606
rect 9254 11578 9282 11583
rect 9254 11531 9282 11550
rect 9198 11466 9226 11471
rect 9366 11466 9394 11471
rect 9198 11419 9226 11438
rect 9254 11438 9366 11466
rect 9142 11326 9226 11354
rect 9198 11186 9226 11326
rect 9198 11153 9226 11158
rect 9142 11129 9170 11135
rect 9142 11103 9143 11129
rect 9169 11103 9170 11129
rect 9142 11074 9170 11103
rect 9198 11074 9226 11079
rect 9142 11046 9198 11074
rect 9198 11041 9226 11046
rect 9198 10794 9226 10799
rect 9254 10794 9282 11438
rect 9366 11433 9394 11438
rect 9310 11242 9338 11247
rect 9310 11129 9338 11214
rect 9310 11103 9311 11129
rect 9337 11103 9338 11129
rect 9310 11097 9338 11103
rect 9534 11073 9562 11830
rect 9590 11857 9618 11863
rect 9590 11831 9591 11857
rect 9617 11831 9618 11857
rect 9590 11746 9618 11831
rect 9590 11713 9618 11718
rect 9702 11857 9730 11863
rect 9702 11831 9703 11857
rect 9729 11831 9730 11857
rect 9534 11047 9535 11073
rect 9561 11047 9562 11073
rect 9534 11018 9562 11047
rect 9534 10985 9562 10990
rect 9702 11690 9730 11831
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9310 10962 9338 10967
rect 9310 10905 9338 10934
rect 9310 10879 9311 10905
rect 9337 10879 9338 10905
rect 9310 10873 9338 10879
rect 9198 10793 9282 10794
rect 9198 10767 9199 10793
rect 9225 10767 9282 10793
rect 9198 10766 9282 10767
rect 9198 10761 9226 10766
rect 9086 10374 9170 10402
rect 9086 10066 9114 10071
rect 9086 10019 9114 10038
rect 9142 9954 9170 10374
rect 9254 10066 9282 10766
rect 9254 10033 9282 10038
rect 9422 10850 9450 10855
rect 9422 10009 9450 10822
rect 9534 10794 9562 10799
rect 9534 10747 9562 10766
rect 9702 10626 9730 11662
rect 9926 11578 9954 11583
rect 9926 11531 9954 11550
rect 10318 11578 10346 12278
rect 10430 12273 10458 12278
rect 9870 11466 9898 11471
rect 9870 11419 9898 11438
rect 9758 11186 9786 11191
rect 9758 11129 9786 11158
rect 10038 11186 10066 11191
rect 10262 11186 10290 11205
rect 10038 11185 10178 11186
rect 10038 11159 10039 11185
rect 10065 11159 10178 11185
rect 10038 11158 10178 11159
rect 10038 11153 10066 11158
rect 9758 11103 9759 11129
rect 9785 11103 9786 11129
rect 9758 10962 9786 11103
rect 9870 11130 9898 11135
rect 9870 11083 9898 11102
rect 10094 11074 10122 11079
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9758 10929 9786 10934
rect 9758 10794 9786 10799
rect 9758 10747 9786 10766
rect 10038 10794 10066 10799
rect 9702 10598 9786 10626
rect 9422 9983 9423 10009
rect 9449 9983 9450 10009
rect 9422 9977 9450 9983
rect 9590 10066 9618 10071
rect 9590 10009 9618 10038
rect 9590 9983 9591 10009
rect 9617 9983 9618 10009
rect 9142 9907 9170 9926
rect 9478 9954 9506 9959
rect 9030 9809 9058 9814
rect 9198 9898 9226 9903
rect 8806 9591 8807 9617
rect 8833 9591 8834 9617
rect 8806 9585 8834 9591
rect 9030 9618 9058 9623
rect 8974 9505 9002 9511
rect 8974 9479 8975 9505
rect 9001 9479 9002 9505
rect 8694 8890 8722 8895
rect 8694 8843 8722 8862
rect 8750 8441 8778 8447
rect 8750 8415 8751 8441
rect 8777 8415 8778 8441
rect 8750 8386 8778 8415
rect 8750 8353 8778 8358
rect 8414 8049 8498 8050
rect 8414 8023 8415 8049
rect 8441 8023 8498 8049
rect 8414 8022 8498 8023
rect 8750 8049 8778 8055
rect 8750 8023 8751 8049
rect 8777 8023 8778 8049
rect 8414 8017 8442 8022
rect 7854 7961 7882 7966
rect 8526 7994 8554 7999
rect 8526 7947 8554 7966
rect 8470 7937 8498 7943
rect 8470 7911 8471 7937
rect 8497 7911 8498 7937
rect 7462 7611 7490 7630
rect 7854 7658 7882 7663
rect 6062 7602 6090 7607
rect 6006 7601 6090 7602
rect 6006 7575 6063 7601
rect 6089 7575 6090 7601
rect 6006 7574 6090 7575
rect 6062 7569 6090 7574
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7854 7265 7882 7630
rect 8470 7574 8498 7911
rect 8750 7769 8778 8023
rect 8750 7743 8751 7769
rect 8777 7743 8778 7769
rect 8750 7737 8778 7743
rect 8190 7546 8498 7574
rect 8862 7713 8890 7719
rect 8862 7687 8863 7713
rect 8889 7687 8890 7713
rect 8190 7321 8218 7546
rect 8190 7295 8191 7321
rect 8217 7295 8218 7321
rect 8190 7289 8218 7295
rect 8862 7322 8890 7687
rect 8918 7714 8946 7719
rect 8974 7714 9002 9479
rect 9030 8833 9058 9590
rect 9198 9561 9226 9870
rect 9198 9535 9199 9561
rect 9225 9535 9226 9561
rect 9198 9529 9226 9535
rect 9366 9673 9394 9679
rect 9366 9647 9367 9673
rect 9393 9647 9394 9673
rect 9254 9226 9282 9231
rect 9254 9179 9282 9198
rect 9366 9226 9394 9647
rect 9422 9618 9450 9623
rect 9478 9618 9506 9926
rect 9422 9617 9506 9618
rect 9422 9591 9423 9617
rect 9449 9591 9506 9617
rect 9422 9590 9506 9591
rect 9534 9897 9562 9903
rect 9534 9871 9535 9897
rect 9561 9871 9562 9897
rect 9422 9585 9450 9590
rect 9422 9226 9450 9231
rect 9366 9225 9450 9226
rect 9366 9199 9423 9225
rect 9449 9199 9450 9225
rect 9366 9198 9450 9199
rect 9030 8807 9031 8833
rect 9057 8807 9058 8833
rect 9030 8386 9058 8807
rect 9366 8833 9394 9198
rect 9422 9193 9450 9198
rect 9534 9114 9562 9871
rect 9590 9617 9618 9983
rect 9590 9591 9591 9617
rect 9617 9591 9618 9617
rect 9590 9585 9618 9591
rect 9702 10010 9730 10015
rect 9646 9226 9674 9231
rect 9702 9226 9730 9982
rect 9758 9506 9786 10598
rect 10038 10401 10066 10766
rect 10038 10375 10039 10401
rect 10065 10375 10066 10401
rect 10038 10369 10066 10375
rect 10094 10402 10122 11046
rect 10094 10369 10122 10374
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10150 10178 10178 11158
rect 10262 11153 10290 11158
rect 9918 10173 10050 10178
rect 10094 10150 10178 10178
rect 10262 11074 10290 11079
rect 10318 11074 10346 11550
rect 10290 11046 10346 11074
rect 10374 11690 10402 11695
rect 10374 11129 10402 11662
rect 10486 11634 10514 11639
rect 10486 11587 10514 11606
rect 10374 11103 10375 11129
rect 10401 11103 10402 11129
rect 10094 10122 10122 10150
rect 10038 10094 10122 10122
rect 10262 10121 10290 11046
rect 10374 11018 10402 11103
rect 10374 10985 10402 10990
rect 10598 11577 10626 11583
rect 10598 11551 10599 11577
rect 10625 11551 10626 11577
rect 10262 10095 10263 10121
rect 10289 10095 10290 10121
rect 9870 9954 9898 9959
rect 9870 9907 9898 9926
rect 10038 9618 10066 10094
rect 10262 10089 10290 10095
rect 10374 10402 10402 10407
rect 10374 10065 10402 10374
rect 10374 10039 10375 10065
rect 10401 10039 10402 10065
rect 10374 10033 10402 10039
rect 10318 10010 10346 10015
rect 10318 9963 10346 9982
rect 10598 9954 10626 11551
rect 10710 11298 10738 12614
rect 10766 12609 10794 12614
rect 10710 11265 10738 11270
rect 10766 11578 10794 11583
rect 10766 11242 10794 11550
rect 10822 11521 10850 12670
rect 10878 12665 10906 12670
rect 10990 12698 11018 12703
rect 11046 12698 11074 13174
rect 11102 12698 11130 12703
rect 11046 12697 11130 12698
rect 11046 12671 11103 12697
rect 11129 12671 11130 12697
rect 11046 12670 11130 12671
rect 10990 12651 11018 12670
rect 11102 12665 11130 12670
rect 11158 12697 11186 13286
rect 11158 12671 11159 12697
rect 11185 12671 11186 12697
rect 11158 12586 11186 12671
rect 11158 12553 11186 12558
rect 11270 13202 11298 13207
rect 11270 13145 11298 13174
rect 11270 13119 11271 13145
rect 11297 13119 11298 13145
rect 11270 11969 11298 13119
rect 11438 13034 11466 13454
rect 11550 13257 11578 13903
rect 11718 13929 11746 13935
rect 11718 13903 11719 13929
rect 11745 13903 11746 13929
rect 11718 13482 11746 13903
rect 12110 13593 12138 14014
rect 12110 13567 12111 13593
rect 12137 13567 12138 13593
rect 12110 13561 12138 13567
rect 11718 13449 11746 13454
rect 11550 13231 11551 13257
rect 11577 13231 11578 13257
rect 11550 13225 11578 13231
rect 12334 13425 12362 13431
rect 12334 13399 12335 13425
rect 12361 13399 12362 13425
rect 11830 13202 11858 13207
rect 12334 13202 12362 13399
rect 11858 13174 11970 13202
rect 11830 13155 11858 13174
rect 11494 13146 11522 13151
rect 11494 13099 11522 13118
rect 11550 13034 11578 13039
rect 11438 13033 11578 13034
rect 11438 13007 11551 13033
rect 11577 13007 11578 13033
rect 11438 13006 11578 13007
rect 11550 13001 11578 13006
rect 11942 12753 11970 13174
rect 12334 13169 12362 13174
rect 12950 13202 12978 13207
rect 11942 12727 11943 12753
rect 11969 12727 11970 12753
rect 11942 12721 11970 12727
rect 12166 13090 12194 13095
rect 12166 12473 12194 13062
rect 12670 13090 12698 13095
rect 12670 13043 12698 13062
rect 12614 13034 12642 13039
rect 12334 13033 12642 13034
rect 12334 13007 12615 13033
rect 12641 13007 12642 13033
rect 12334 13006 12642 13007
rect 12334 12809 12362 13006
rect 12614 13001 12642 13006
rect 12334 12783 12335 12809
rect 12361 12783 12362 12809
rect 12334 12777 12362 12783
rect 12950 12642 12978 13174
rect 13398 12810 13426 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 20118 18129 20146 18135
rect 20118 18103 20119 18129
rect 20145 18103 20146 18129
rect 20118 17850 20146 18103
rect 20118 17817 20146 17822
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 20118 13425 20146 13431
rect 20118 13399 20119 13425
rect 20145 13399 20146 13425
rect 20118 13146 20146 13399
rect 20118 13113 20146 13118
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 12278 12586 12306 12591
rect 12166 12447 12167 12473
rect 12193 12447 12194 12473
rect 12166 12441 12194 12447
rect 12222 12474 12250 12479
rect 12222 12427 12250 12446
rect 12278 12473 12306 12558
rect 12278 12447 12279 12473
rect 12305 12447 12306 12473
rect 12278 12441 12306 12447
rect 11998 12362 12026 12367
rect 11270 11943 11271 11969
rect 11297 11943 11298 11969
rect 11270 11937 11298 11943
rect 11718 12361 12026 12362
rect 11718 12335 11999 12361
rect 12025 12335 12026 12361
rect 11718 12334 12026 12335
rect 11662 11913 11690 11919
rect 11662 11887 11663 11913
rect 11689 11887 11690 11913
rect 11158 11802 11186 11807
rect 10878 11690 10906 11695
rect 10878 11643 10906 11662
rect 11158 11689 11186 11774
rect 11158 11663 11159 11689
rect 11185 11663 11186 11689
rect 11158 11657 11186 11663
rect 10822 11495 10823 11521
rect 10849 11495 10850 11521
rect 10822 11489 10850 11495
rect 11046 11577 11074 11583
rect 11046 11551 11047 11577
rect 11073 11551 11074 11577
rect 10766 11209 10794 11214
rect 10990 11298 11018 11303
rect 10710 11074 10738 11079
rect 10710 11027 10738 11046
rect 10878 11073 10906 11079
rect 10878 11047 10879 11073
rect 10905 11047 10906 11073
rect 10878 10962 10906 11047
rect 10766 10402 10794 10407
rect 10878 10402 10906 10934
rect 10766 10401 10906 10402
rect 10766 10375 10767 10401
rect 10793 10375 10906 10401
rect 10766 10374 10906 10375
rect 10934 10402 10962 10407
rect 10766 10369 10794 10374
rect 10934 10355 10962 10374
rect 10710 10290 10738 10295
rect 10710 10243 10738 10262
rect 10990 10121 11018 11270
rect 11046 11186 11074 11551
rect 11606 11578 11634 11583
rect 11214 11466 11242 11471
rect 11046 11153 11074 11158
rect 11158 11465 11242 11466
rect 11158 11439 11215 11465
rect 11241 11439 11242 11465
rect 11158 11438 11242 11439
rect 11102 11074 11130 11079
rect 11158 11074 11186 11438
rect 11214 11433 11242 11438
rect 11130 11046 11186 11074
rect 11214 11185 11242 11191
rect 11494 11186 11522 11191
rect 11214 11159 11215 11185
rect 11241 11159 11242 11185
rect 11102 11027 11130 11046
rect 11214 10850 11242 11159
rect 11214 10817 11242 10822
rect 11438 11185 11522 11186
rect 11438 11159 11495 11185
rect 11521 11159 11522 11185
rect 11438 11158 11522 11159
rect 11382 10402 11410 10407
rect 11382 10355 11410 10374
rect 11158 10346 11186 10351
rect 11158 10299 11186 10318
rect 11438 10345 11466 11158
rect 11494 11153 11522 11158
rect 11438 10319 11439 10345
rect 11465 10319 11466 10345
rect 10990 10095 10991 10121
rect 11017 10095 11018 10121
rect 10626 9926 10738 9954
rect 10598 9921 10626 9926
rect 10038 9571 10066 9590
rect 9870 9506 9898 9511
rect 9758 9505 9898 9506
rect 9758 9479 9871 9505
rect 9897 9479 9898 9505
rect 9758 9478 9898 9479
rect 9758 9281 9786 9478
rect 9870 9473 9898 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9814 9338 9842 9343
rect 9814 9291 9842 9310
rect 10150 9338 10178 9343
rect 9758 9255 9759 9281
rect 9785 9255 9786 9281
rect 9758 9249 9786 9255
rect 10150 9281 10178 9310
rect 10150 9255 10151 9281
rect 10177 9255 10178 9281
rect 10150 9249 10178 9255
rect 9646 9225 9730 9226
rect 9646 9199 9647 9225
rect 9673 9199 9730 9225
rect 9646 9198 9730 9199
rect 10038 9226 10066 9231
rect 9646 9193 9674 9198
rect 9982 9114 10010 9119
rect 9562 9086 9618 9114
rect 9534 9067 9562 9086
rect 9590 9058 9618 9086
rect 9870 9086 9982 9114
rect 9590 9030 9674 9058
rect 9366 8807 9367 8833
rect 9393 8807 9394 8833
rect 9366 8554 9394 8807
rect 9646 8833 9674 9030
rect 9870 8945 9898 9086
rect 9982 9067 10010 9086
rect 9870 8919 9871 8945
rect 9897 8919 9898 8945
rect 9870 8913 9898 8919
rect 9926 8946 9954 8951
rect 10038 8946 10066 9198
rect 10318 9225 10346 9231
rect 10318 9199 10319 9225
rect 10345 9199 10346 9225
rect 10318 9170 10346 9199
rect 9926 8945 10066 8946
rect 9926 8919 9927 8945
rect 9953 8919 10066 8945
rect 9926 8918 10066 8919
rect 10206 9142 10318 9170
rect 9926 8913 9954 8918
rect 10206 8890 10234 9142
rect 10318 9137 10346 9142
rect 10374 9225 10402 9231
rect 10374 9199 10375 9225
rect 10401 9199 10402 9225
rect 9646 8807 9647 8833
rect 9673 8807 9674 8833
rect 9646 8801 9674 8807
rect 10094 8862 10234 8890
rect 9590 8778 9618 8783
rect 9590 8731 9618 8750
rect 10038 8777 10066 8783
rect 10038 8751 10039 8777
rect 10065 8751 10066 8777
rect 9534 8722 9562 8727
rect 9534 8675 9562 8694
rect 10038 8722 10066 8751
rect 10038 8689 10066 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9366 8521 9394 8526
rect 9086 8498 9114 8503
rect 9086 8451 9114 8470
rect 9058 8358 9114 8386
rect 9030 8353 9058 8358
rect 8946 7686 9002 7714
rect 9086 8050 9114 8358
rect 8918 7667 8946 7686
rect 9086 7657 9114 8022
rect 10094 7993 10122 8862
rect 10206 8833 10234 8862
rect 10374 8890 10402 9199
rect 10374 8857 10402 8862
rect 10430 9225 10458 9231
rect 10430 9199 10431 9225
rect 10457 9199 10458 9225
rect 10430 9058 10458 9199
rect 10206 8807 10207 8833
rect 10233 8807 10234 8833
rect 10206 8801 10234 8807
rect 10150 8778 10178 8783
rect 10150 8386 10178 8750
rect 10318 8778 10346 8783
rect 10430 8778 10458 9030
rect 10710 8889 10738 9926
rect 10934 9730 10962 9735
rect 10878 9281 10906 9287
rect 10878 9255 10879 9281
rect 10905 9255 10906 9281
rect 10710 8863 10711 8889
rect 10737 8863 10738 8889
rect 10710 8857 10738 8863
rect 10766 9225 10794 9231
rect 10766 9199 10767 9225
rect 10793 9199 10794 9225
rect 10318 8777 10458 8778
rect 10318 8751 10319 8777
rect 10345 8751 10458 8777
rect 10318 8750 10458 8751
rect 10318 8745 10346 8750
rect 10262 8721 10290 8727
rect 10262 8695 10263 8721
rect 10289 8695 10290 8721
rect 10262 8498 10290 8695
rect 10262 8465 10290 8470
rect 10542 8442 10570 8447
rect 10150 8385 10234 8386
rect 10150 8359 10151 8385
rect 10177 8359 10234 8385
rect 10150 8358 10234 8359
rect 10150 8353 10178 8358
rect 10150 8050 10178 8055
rect 10150 8003 10178 8022
rect 10094 7967 10095 7993
rect 10121 7967 10122 7993
rect 10094 7961 10122 7967
rect 9982 7938 10010 7943
rect 9478 7937 10010 7938
rect 9478 7911 9983 7937
rect 10009 7911 10010 7937
rect 9478 7910 10010 7911
rect 9478 7713 9506 7910
rect 9982 7905 10010 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9478 7687 9479 7713
rect 9505 7687 9506 7713
rect 9478 7681 9506 7687
rect 9086 7631 9087 7657
rect 9113 7631 9114 7657
rect 9086 7625 9114 7631
rect 7854 7239 7855 7265
rect 7881 7239 7882 7265
rect 7854 7233 7882 7239
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8862 4214 8890 7294
rect 9254 7322 9282 7327
rect 9254 7275 9282 7294
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 8806 4186 8890 4214
rect 10206 4214 10234 8358
rect 10542 7601 10570 8414
rect 10766 8050 10794 9199
rect 10878 8834 10906 9255
rect 10934 9281 10962 9702
rect 10934 9255 10935 9281
rect 10961 9255 10962 9281
rect 10934 9249 10962 9255
rect 10990 9226 11018 10095
rect 11102 10122 11130 10127
rect 11102 10075 11130 10094
rect 11438 10122 11466 10319
rect 11158 10066 11186 10071
rect 11158 10019 11186 10038
rect 11214 9730 11242 9735
rect 11214 9683 11242 9702
rect 10990 9193 11018 9198
rect 11102 9618 11130 9623
rect 11102 9058 11130 9590
rect 11270 9562 11298 9567
rect 11438 9562 11466 10094
rect 11606 9618 11634 11550
rect 11662 11521 11690 11887
rect 11718 11802 11746 12334
rect 11998 12329 12026 12334
rect 12110 12361 12138 12367
rect 12110 12335 12111 12361
rect 12137 12335 12138 12361
rect 11718 11689 11746 11774
rect 11718 11663 11719 11689
rect 11745 11663 11746 11689
rect 11718 11657 11746 11663
rect 11662 11495 11663 11521
rect 11689 11495 11690 11521
rect 11662 11489 11690 11495
rect 11886 11634 11914 11639
rect 11830 11465 11858 11471
rect 11830 11439 11831 11465
rect 11857 11439 11858 11465
rect 11774 11186 11802 11191
rect 11718 11185 11802 11186
rect 11718 11159 11775 11185
rect 11801 11159 11802 11185
rect 11718 11158 11802 11159
rect 11662 11129 11690 11135
rect 11662 11103 11663 11129
rect 11689 11103 11690 11129
rect 11662 10066 11690 11103
rect 11718 10962 11746 11158
rect 11774 11153 11802 11158
rect 11774 11074 11802 11079
rect 11830 11074 11858 11439
rect 11886 11241 11914 11606
rect 11886 11215 11887 11241
rect 11913 11215 11914 11241
rect 11886 11209 11914 11215
rect 11942 11578 11970 11583
rect 11774 11073 11858 11074
rect 11774 11047 11775 11073
rect 11801 11047 11858 11073
rect 11774 11046 11858 11047
rect 11774 11041 11802 11046
rect 11886 10962 11914 10967
rect 11718 10934 11802 10962
rect 11718 10794 11746 10799
rect 11718 10737 11746 10766
rect 11718 10711 11719 10737
rect 11745 10711 11746 10737
rect 11718 10705 11746 10711
rect 11774 10457 11802 10934
rect 11774 10431 11775 10457
rect 11801 10431 11802 10457
rect 11774 10425 11802 10431
rect 11886 10401 11914 10934
rect 11886 10375 11887 10401
rect 11913 10375 11914 10401
rect 11886 10369 11914 10375
rect 11662 10033 11690 10038
rect 11718 10346 11746 10351
rect 11662 9618 11690 9623
rect 11606 9617 11690 9618
rect 11606 9591 11663 9617
rect 11689 9591 11690 9617
rect 11606 9590 11690 9591
rect 11662 9585 11690 9590
rect 11270 9561 11354 9562
rect 11270 9535 11271 9561
rect 11297 9535 11354 9561
rect 11270 9534 11354 9535
rect 11438 9534 11634 9562
rect 11270 9529 11298 9534
rect 11270 9338 11298 9343
rect 11158 9310 11270 9338
rect 11158 9169 11186 9310
rect 11270 9305 11298 9310
rect 11326 9226 11354 9534
rect 11550 9282 11578 9287
rect 11494 9254 11550 9282
rect 11326 9225 11466 9226
rect 11326 9199 11327 9225
rect 11353 9199 11466 9225
rect 11326 9198 11466 9199
rect 11326 9193 11354 9198
rect 11158 9143 11159 9169
rect 11185 9143 11186 9169
rect 11158 9137 11186 9143
rect 11102 9030 11298 9058
rect 11046 8946 11074 8951
rect 10878 8787 10906 8806
rect 10934 8889 10962 8895
rect 10934 8863 10935 8889
rect 10961 8863 10962 8889
rect 10878 8442 10906 8447
rect 10934 8442 10962 8863
rect 11046 8553 11074 8918
rect 11270 8945 11298 9030
rect 11270 8919 11271 8945
rect 11297 8919 11298 8945
rect 11270 8913 11298 8919
rect 11438 8946 11466 9198
rect 11438 8899 11466 8918
rect 11046 8527 11047 8553
rect 11073 8527 11074 8553
rect 11046 8521 11074 8527
rect 11382 8834 11410 8839
rect 11382 8497 11410 8806
rect 11494 8722 11522 9254
rect 11550 9235 11578 9254
rect 11382 8471 11383 8497
rect 11409 8471 11410 8497
rect 11382 8465 11410 8471
rect 11438 8694 11522 8722
rect 11550 8834 11578 8839
rect 10906 8414 10962 8442
rect 10878 8395 10906 8414
rect 10766 8017 10794 8022
rect 11438 8329 11466 8694
rect 11438 8303 11439 8329
rect 11465 8303 11466 8329
rect 11102 7714 11130 7719
rect 11438 7714 11466 8303
rect 11494 7994 11522 7999
rect 11550 7994 11578 8806
rect 11606 8498 11634 9534
rect 11718 9338 11746 10318
rect 11942 10121 11970 11550
rect 12110 11578 12138 12335
rect 12726 12026 12754 12031
rect 12110 11545 12138 11550
rect 12614 12025 12754 12026
rect 12614 11999 12727 12025
rect 12753 11999 12754 12025
rect 12614 11998 12754 11999
rect 12614 11690 12642 11998
rect 12726 11993 12754 11998
rect 12950 12025 12978 12614
rect 13342 12809 13426 12810
rect 13342 12783 13399 12809
rect 13425 12783 13426 12809
rect 13342 12782 13426 12783
rect 13342 12474 13370 12782
rect 13398 12777 13426 12782
rect 13342 12441 13370 12446
rect 13398 12642 13426 12647
rect 13622 12642 13650 12647
rect 13426 12641 13650 12642
rect 13426 12615 13623 12641
rect 13649 12615 13650 12641
rect 13426 12614 13650 12615
rect 12950 11999 12951 12025
rect 12977 11999 12978 12025
rect 12950 11993 12978 11999
rect 11998 11186 12026 11191
rect 11998 11139 12026 11158
rect 12278 11185 12306 11191
rect 12278 11159 12279 11185
rect 12305 11159 12306 11185
rect 12166 11130 12194 11135
rect 12166 11074 12194 11102
rect 12110 11073 12194 11074
rect 12110 11047 12167 11073
rect 12193 11047 12194 11073
rect 12110 11046 12194 11047
rect 11942 10095 11943 10121
rect 11969 10095 11970 10121
rect 11942 10089 11970 10095
rect 11998 10346 12026 10351
rect 11886 10065 11914 10071
rect 11886 10039 11887 10065
rect 11913 10039 11914 10065
rect 11774 9506 11802 9511
rect 11774 9505 11858 9506
rect 11774 9479 11775 9505
rect 11801 9479 11858 9505
rect 11774 9478 11858 9479
rect 11774 9473 11802 9478
rect 11718 9225 11746 9310
rect 11718 9199 11719 9225
rect 11745 9199 11746 9225
rect 11718 9193 11746 9199
rect 11830 9114 11858 9478
rect 11886 9505 11914 10039
rect 11998 10065 12026 10318
rect 11998 10039 11999 10065
rect 12025 10039 12026 10065
rect 11998 10033 12026 10039
rect 11942 9730 11970 9735
rect 11942 9683 11970 9702
rect 11886 9479 11887 9505
rect 11913 9479 11914 9505
rect 11886 9282 11914 9479
rect 11886 9249 11914 9254
rect 11718 8946 11746 8951
rect 11718 8833 11746 8918
rect 11718 8807 11719 8833
rect 11745 8807 11746 8833
rect 11718 8801 11746 8807
rect 11830 8722 11858 9086
rect 11886 9170 11914 9175
rect 11886 8834 11914 9142
rect 12054 9058 12082 9063
rect 12110 9058 12138 11046
rect 12166 11041 12194 11046
rect 12278 10962 12306 11159
rect 12614 11186 12642 11662
rect 12726 11914 12754 11919
rect 12726 11689 12754 11886
rect 12726 11663 12727 11689
rect 12753 11663 12754 11689
rect 12726 11657 12754 11663
rect 12670 11634 12698 11639
rect 12670 11587 12698 11606
rect 12950 11634 12978 11639
rect 12950 11587 12978 11606
rect 12782 11578 12810 11583
rect 12782 11531 12810 11550
rect 13230 11578 13258 11583
rect 13342 11578 13370 11583
rect 13398 11578 13426 12614
rect 13622 12609 13650 12614
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 18942 11969 18970 11975
rect 18942 11943 18943 11969
rect 18969 11943 18970 11969
rect 13566 11914 13594 11919
rect 13566 11867 13594 11886
rect 13622 11857 13650 11863
rect 13622 11831 13623 11857
rect 13649 11831 13650 11857
rect 13258 11550 13314 11578
rect 13230 11545 13258 11550
rect 12614 11153 12642 11158
rect 13062 11465 13090 11471
rect 13062 11439 13063 11465
rect 13089 11439 13090 11465
rect 12726 11074 12754 11079
rect 12670 10962 12698 10967
rect 12306 10934 12418 10962
rect 12278 10929 12306 10934
rect 12166 10850 12194 10855
rect 12166 10402 12194 10822
rect 12166 10345 12194 10374
rect 12390 10401 12418 10934
rect 12614 10794 12642 10799
rect 12614 10747 12642 10766
rect 12670 10682 12698 10934
rect 12614 10654 12698 10682
rect 12614 10457 12642 10654
rect 12726 10458 12754 11046
rect 12614 10431 12615 10457
rect 12641 10431 12642 10457
rect 12614 10425 12642 10431
rect 12670 10430 12754 10458
rect 12894 11018 12922 11023
rect 12390 10375 12391 10401
rect 12417 10375 12418 10401
rect 12390 10369 12418 10375
rect 12166 10319 12167 10345
rect 12193 10319 12194 10345
rect 12166 10313 12194 10319
rect 12502 10346 12530 10351
rect 12502 10299 12530 10318
rect 12670 10345 12698 10430
rect 12838 10402 12866 10407
rect 12838 10355 12866 10374
rect 12670 10319 12671 10345
rect 12697 10319 12698 10345
rect 12670 10313 12698 10319
rect 12726 10346 12754 10351
rect 12726 10093 12754 10318
rect 12670 10065 12698 10071
rect 12670 10039 12671 10065
rect 12697 10039 12698 10065
rect 12726 10067 12727 10093
rect 12753 10067 12754 10093
rect 12726 10061 12754 10067
rect 12894 10065 12922 10990
rect 13062 10962 13090 11439
rect 13118 11466 13146 11471
rect 13118 11419 13146 11438
rect 13174 11185 13202 11191
rect 13174 11159 13175 11185
rect 13201 11159 13202 11185
rect 13174 11130 13202 11159
rect 13286 11186 13314 11550
rect 13342 11577 13398 11578
rect 13342 11551 13343 11577
rect 13369 11551 13398 11577
rect 13342 11550 13398 11551
rect 13342 11545 13370 11550
rect 13398 11531 13426 11550
rect 13454 11634 13482 11639
rect 13622 11634 13650 11831
rect 13678 11634 13706 11639
rect 13622 11633 13706 11634
rect 13622 11607 13679 11633
rect 13705 11607 13706 11633
rect 13622 11606 13706 11607
rect 13342 11186 13370 11191
rect 13286 11185 13370 11186
rect 13286 11159 13343 11185
rect 13369 11159 13370 11185
rect 13286 11158 13370 11159
rect 13342 11153 13370 11158
rect 13174 11097 13202 11102
rect 13454 11129 13482 11606
rect 13678 11601 13706 11606
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 14742 11521 14770 11527
rect 14742 11495 14743 11521
rect 14769 11495 14770 11521
rect 14742 11466 14770 11495
rect 14966 11522 14994 11527
rect 14994 11494 15050 11522
rect 14966 11475 14994 11494
rect 14742 11433 14770 11438
rect 13454 11103 13455 11129
rect 13481 11103 13482 11129
rect 13062 10929 13090 10934
rect 13286 11073 13314 11079
rect 13286 11047 13287 11073
rect 13313 11047 13314 11073
rect 13286 10570 13314 11047
rect 13286 10537 13314 10542
rect 13006 10346 13034 10351
rect 13006 10299 13034 10318
rect 13454 10346 13482 11103
rect 13622 11185 13650 11191
rect 13622 11159 13623 11185
rect 13649 11159 13650 11185
rect 13622 10962 13650 11159
rect 13678 11186 13706 11191
rect 14238 11186 14266 11191
rect 13678 11185 14266 11186
rect 13678 11159 13679 11185
rect 13705 11159 14239 11185
rect 14265 11159 14266 11185
rect 13678 11158 14266 11159
rect 13678 11153 13706 11158
rect 14238 11153 14266 11158
rect 14294 11130 14322 11135
rect 14294 11083 14322 11102
rect 14798 11130 14826 11135
rect 13622 10929 13650 10934
rect 14686 11018 14714 11023
rect 13734 10570 13762 10575
rect 13566 10402 13594 10407
rect 13510 10346 13538 10351
rect 13482 10345 13538 10346
rect 13482 10319 13511 10345
rect 13537 10319 13538 10345
rect 13482 10318 13538 10319
rect 13454 10299 13482 10318
rect 13510 10313 13538 10318
rect 13566 10345 13594 10374
rect 13566 10319 13567 10345
rect 13593 10319 13594 10345
rect 13566 10313 13594 10319
rect 12670 10010 12698 10039
rect 12894 10039 12895 10065
rect 12921 10039 12922 10065
rect 12670 9982 12754 10010
rect 12726 9954 12754 9982
rect 12894 9954 12922 10039
rect 13230 10290 13258 10295
rect 12726 9926 12922 9954
rect 13006 10009 13034 10015
rect 13006 9983 13007 10009
rect 13033 9983 13034 10009
rect 12082 9030 12138 9058
rect 12670 9897 12698 9903
rect 12670 9871 12671 9897
rect 12697 9871 12698 9897
rect 12054 9025 12082 9030
rect 11886 8801 11914 8806
rect 11886 8722 11914 8727
rect 11830 8694 11886 8722
rect 11886 8675 11914 8694
rect 12614 8554 12642 8559
rect 12558 8553 12642 8554
rect 12558 8527 12615 8553
rect 12641 8527 12642 8553
rect 12558 8526 12642 8527
rect 11830 8498 11858 8503
rect 11606 8470 11830 8498
rect 11662 8050 11690 8055
rect 11662 8003 11690 8022
rect 11494 7993 11578 7994
rect 11494 7967 11495 7993
rect 11521 7967 11578 7993
rect 11494 7966 11578 7967
rect 11830 7993 11858 8470
rect 12558 8105 12586 8526
rect 12614 8521 12642 8526
rect 12670 8554 12698 9871
rect 13006 9730 13034 9983
rect 13230 10009 13258 10262
rect 13678 10290 13706 10295
rect 13678 10243 13706 10262
rect 13734 10065 13762 10542
rect 13734 10039 13735 10065
rect 13761 10039 13762 10065
rect 13734 10033 13762 10039
rect 14294 10402 14322 10407
rect 13230 9983 13231 10009
rect 13257 9983 13258 10009
rect 13230 9977 13258 9983
rect 13342 10009 13370 10015
rect 13342 9983 13343 10009
rect 13369 9983 13370 10009
rect 13118 9953 13146 9959
rect 13118 9927 13119 9953
rect 13145 9927 13146 9953
rect 13118 9730 13146 9927
rect 13118 9702 13258 9730
rect 13006 9697 13034 9702
rect 13230 9673 13258 9702
rect 13230 9647 13231 9673
rect 13257 9647 13258 9673
rect 13230 9641 13258 9647
rect 12894 9617 12922 9623
rect 12894 9591 12895 9617
rect 12921 9591 12922 9617
rect 12894 9226 12922 9591
rect 12894 9193 12922 9198
rect 13286 9226 13314 9231
rect 13342 9226 13370 9983
rect 14294 9673 14322 10374
rect 14294 9647 14295 9673
rect 14321 9647 14322 9673
rect 14294 9641 14322 9647
rect 14574 9618 14602 9623
rect 14574 9571 14602 9590
rect 14686 9617 14714 10990
rect 14798 9953 14826 11102
rect 14798 9927 14799 9953
rect 14825 9927 14826 9953
rect 14798 9921 14826 9927
rect 15022 10737 15050 11494
rect 18942 11466 18970 11943
rect 20006 11802 20034 11999
rect 20006 11769 20034 11774
rect 18942 11433 18970 11438
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 15022 10711 15023 10737
rect 15049 10711 15050 10737
rect 15022 9953 15050 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 18830 10402 18858 10407
rect 18830 10355 18858 10374
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 15022 9927 15023 9953
rect 15049 9927 15050 9953
rect 14686 9591 14687 9617
rect 14713 9591 14714 9617
rect 14686 9585 14714 9591
rect 13314 9198 13370 9226
rect 13622 9506 13650 9511
rect 13622 9225 13650 9478
rect 14630 9506 14658 9511
rect 14630 9459 14658 9478
rect 14798 9505 14826 9511
rect 14798 9479 14799 9505
rect 14825 9479 14826 9505
rect 13622 9199 13623 9225
rect 13649 9199 13650 9225
rect 13230 8834 13258 8839
rect 12670 8441 12698 8526
rect 12782 8722 12810 8727
rect 12670 8415 12671 8441
rect 12697 8415 12698 8441
rect 12670 8409 12698 8415
rect 12726 8442 12754 8447
rect 12558 8079 12559 8105
rect 12585 8079 12586 8105
rect 12558 8073 12586 8079
rect 11998 8050 12026 8055
rect 12026 8022 12194 8050
rect 11998 8003 12026 8022
rect 11830 7967 11831 7993
rect 11857 7967 11858 7993
rect 11494 7961 11522 7966
rect 11830 7961 11858 7967
rect 11102 7713 11466 7714
rect 11102 7687 11103 7713
rect 11129 7687 11466 7713
rect 11102 7686 11466 7687
rect 11102 7681 11130 7686
rect 10766 7658 10794 7663
rect 10766 7611 10794 7630
rect 10542 7575 10543 7601
rect 10569 7575 10570 7601
rect 10542 7569 10570 7575
rect 12166 7601 12194 8022
rect 12166 7575 12167 7601
rect 12193 7575 12194 7601
rect 12166 7569 12194 7575
rect 12222 8049 12250 8055
rect 12222 8023 12223 8049
rect 12249 8023 12250 8049
rect 12222 7658 12250 8023
rect 12222 7574 12250 7630
rect 12726 7658 12754 8414
rect 12782 8441 12810 8694
rect 13230 8553 13258 8806
rect 13230 8527 13231 8553
rect 13257 8527 13258 8553
rect 13230 8521 13258 8527
rect 12950 8498 12978 8503
rect 12950 8451 12978 8470
rect 13286 8498 13314 9198
rect 13622 9193 13650 9199
rect 14070 9282 14098 9287
rect 13958 9170 13986 9175
rect 13902 8777 13930 8783
rect 13902 8751 13903 8777
rect 13929 8751 13930 8777
rect 13342 8554 13370 8559
rect 13342 8507 13370 8526
rect 13286 8465 13314 8470
rect 12782 8415 12783 8441
rect 12809 8415 12810 8441
rect 12782 8409 12810 8415
rect 13566 8441 13594 8447
rect 13566 8415 13567 8441
rect 13593 8415 13594 8441
rect 13286 8385 13314 8391
rect 13286 8359 13287 8385
rect 13313 8359 13314 8385
rect 13062 8330 13090 8335
rect 13062 8283 13090 8302
rect 13118 7714 13146 7719
rect 13286 7714 13314 8359
rect 13566 8274 13594 8415
rect 13734 8442 13762 8447
rect 13734 8395 13762 8414
rect 13566 8241 13594 8246
rect 13734 8330 13762 8335
rect 13622 8106 13650 8111
rect 13622 8059 13650 8078
rect 13734 8049 13762 8302
rect 13734 8023 13735 8049
rect 13761 8023 13762 8049
rect 13734 8017 13762 8023
rect 13846 8106 13874 8111
rect 13846 7993 13874 8078
rect 13846 7967 13847 7993
rect 13873 7967 13874 7993
rect 13846 7961 13874 7967
rect 13902 7994 13930 8751
rect 13958 8777 13986 9142
rect 14070 8833 14098 9254
rect 14798 9282 14826 9479
rect 14798 9249 14826 9254
rect 15022 9506 15050 9927
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 15078 9506 15106 9511
rect 15022 9505 15106 9506
rect 15022 9479 15079 9505
rect 15105 9479 15106 9505
rect 15022 9478 15106 9479
rect 14686 9170 14714 9175
rect 14686 9123 14714 9142
rect 14910 9170 14938 9175
rect 15022 9170 15050 9478
rect 15078 9473 15106 9478
rect 18830 9226 18858 9231
rect 18830 9179 18858 9198
rect 14910 9169 15050 9170
rect 14910 9143 14911 9169
rect 14937 9143 15050 9169
rect 14910 9142 15050 9143
rect 14070 8807 14071 8833
rect 14097 8807 14098 8833
rect 14070 8801 14098 8807
rect 13958 8751 13959 8777
rect 13985 8751 13986 8777
rect 13958 8745 13986 8751
rect 14406 8442 14434 8447
rect 13958 8274 13986 8279
rect 13986 8246 14154 8274
rect 13958 8241 13986 8246
rect 14126 8161 14154 8246
rect 14126 8135 14127 8161
rect 14153 8135 14154 8161
rect 14126 8129 14154 8135
rect 14070 7994 14098 7999
rect 13902 7993 14098 7994
rect 13902 7967 13903 7993
rect 13929 7967 14071 7993
rect 14097 7967 14098 7993
rect 13902 7966 14098 7967
rect 13118 7713 13314 7714
rect 13118 7687 13119 7713
rect 13145 7687 13314 7713
rect 13118 7686 13314 7687
rect 13902 7714 13930 7966
rect 14070 7961 14098 7966
rect 14126 7938 14154 7943
rect 14126 7937 14210 7938
rect 14126 7911 14127 7937
rect 14153 7911 14210 7937
rect 14126 7910 14210 7911
rect 14126 7905 14154 7910
rect 13118 7681 13146 7686
rect 13902 7681 13930 7686
rect 12726 7611 12754 7630
rect 14182 7602 14210 7910
rect 14406 7769 14434 8414
rect 14910 8442 14938 9142
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 14910 8409 14938 8414
rect 18830 8441 18858 8447
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 18830 8162 18858 8415
rect 18830 8129 18858 8134
rect 19950 8385 19978 8391
rect 19950 8359 19951 8385
rect 19977 8359 19978 8385
rect 19950 8106 19978 8359
rect 19950 8073 19978 8078
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 14406 7743 14407 7769
rect 14433 7743 14434 7769
rect 14406 7737 14434 7743
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 12222 7546 12362 7574
rect 14182 7555 14210 7574
rect 18830 7602 18858 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18830 7569 18858 7574
rect 12334 7321 12362 7546
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 12334 7295 12335 7321
rect 12361 7295 12362 7321
rect 12334 7289 12362 7295
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 10206 4186 10402 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8806 1777 8834 4186
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 7854 1666 7882 1671
rect 7742 1665 7882 1666
rect 7742 1639 7855 1665
rect 7881 1639 7882 1665
rect 7742 1638 7882 1639
rect 7742 400 7770 1638
rect 7854 1633 7882 1638
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 9758 1834 9786 1839
rect 9758 400 9786 1806
rect 10374 1777 10402 4186
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 10934 1834 10962 1839
rect 10934 1787 10962 1806
rect 10374 1751 10375 1777
rect 10401 1751 10402 1777
rect 10374 1745 10402 1751
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 7728 0 7784 400
rect 9072 0 9128 400
rect 9744 0 9800 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8414 19110 8442 19138
rect 9030 19137 9058 19138
rect 9030 19111 9031 19137
rect 9031 19111 9057 19137
rect 9057 19111 9058 19137
rect 9030 19110 9058 19111
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 11774 19110 11802 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9422 18718 9450 18746
rect 10038 18745 10066 18746
rect 10038 18719 10039 18745
rect 10039 18719 10065 18745
rect 10065 18719 10066 18745
rect 10038 18718 10066 18719
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 6958 13510 6986 13538
rect 2086 13454 2114 13482
rect 966 12249 994 12250
rect 966 12223 967 12249
rect 967 12223 993 12249
rect 993 12223 994 12249
rect 966 12222 994 12223
rect 966 11241 994 11242
rect 966 11215 967 11241
rect 967 11215 993 11241
rect 993 11215 994 11241
rect 966 11214 994 11215
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 8078 13537 8106 13538
rect 8078 13511 8079 13537
rect 8079 13511 8105 13537
rect 8105 13511 8106 13537
rect 8078 13510 8106 13511
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9198 13510 9226 13538
rect 8806 13454 8834 13482
rect 2142 12361 2170 12362
rect 2142 12335 2143 12361
rect 2143 12335 2169 12361
rect 2169 12335 2170 12361
rect 2142 12334 2170 12335
rect 7294 12446 7322 12474
rect 8134 12473 8162 12474
rect 8134 12447 8135 12473
rect 8135 12447 8161 12473
rect 8161 12447 8162 12473
rect 8134 12446 8162 12447
rect 5670 12334 5698 12362
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 6734 12305 6762 12306
rect 6734 12279 6735 12305
rect 6735 12279 6761 12305
rect 6761 12279 6762 12305
rect 6734 12278 6762 12279
rect 5670 11830 5698 11858
rect 7518 12278 7546 12306
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 6846 11270 6874 11298
rect 2142 11185 2170 11186
rect 2142 11159 2143 11185
rect 2143 11159 2169 11185
rect 2169 11159 2170 11185
rect 2142 11158 2170 11159
rect 5446 11158 5474 11186
rect 2086 10766 2114 10794
rect 6958 11185 6986 11186
rect 6958 11159 6959 11185
rect 6959 11159 6985 11185
rect 6985 11159 6986 11185
rect 6958 11158 6986 11159
rect 6454 10710 6482 10738
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 4998 10457 5026 10458
rect 4998 10431 4999 10457
rect 4999 10431 5025 10457
rect 5025 10431 5026 10457
rect 4998 10430 5026 10431
rect 2142 10401 2170 10402
rect 2142 10375 2143 10401
rect 2143 10375 2169 10401
rect 2169 10375 2170 10401
rect 2142 10374 2170 10375
rect 7126 11857 7154 11858
rect 7126 11831 7127 11857
rect 7127 11831 7153 11857
rect 7153 11831 7154 11857
rect 7126 11830 7154 11831
rect 7070 11270 7098 11298
rect 7238 11606 7266 11634
rect 7350 11521 7378 11522
rect 7350 11495 7351 11521
rect 7351 11495 7377 11521
rect 7377 11495 7378 11521
rect 7350 11494 7378 11495
rect 7630 11158 7658 11186
rect 8302 11662 8330 11690
rect 8190 11494 8218 11522
rect 8806 11662 8834 11690
rect 8358 11185 8386 11186
rect 8358 11159 8359 11185
rect 8359 11159 8385 11185
rect 8385 11159 8386 11185
rect 8358 11158 8386 11159
rect 8134 11129 8162 11130
rect 8134 11103 8135 11129
rect 8135 11103 8161 11129
rect 8161 11103 8162 11129
rect 8134 11102 8162 11103
rect 7238 10990 7266 11018
rect 6902 10710 6930 10738
rect 966 10094 994 10122
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 6062 9870 6090 9898
rect 8470 10878 8498 10906
rect 8526 11438 8554 11466
rect 8862 11158 8890 11186
rect 8526 11102 8554 11130
rect 8918 11102 8946 11130
rect 8974 11550 9002 11578
rect 8806 10905 8834 10906
rect 8806 10879 8807 10905
rect 8807 10879 8833 10905
rect 8833 10879 8834 10905
rect 8806 10878 8834 10879
rect 6566 10430 6594 10458
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6678 10065 6706 10066
rect 6678 10039 6679 10065
rect 6679 10039 6705 10065
rect 6705 10039 6706 10065
rect 6678 10038 6706 10039
rect 4998 9673 5026 9674
rect 4998 9647 4999 9673
rect 4999 9647 5025 9673
rect 5025 9647 5026 9673
rect 4998 9646 5026 9647
rect 2142 9617 2170 9618
rect 2142 9591 2143 9617
rect 2143 9591 2169 9617
rect 2169 9591 2170 9617
rect 2142 9590 2170 9591
rect 966 9422 994 9450
rect 5838 9310 5866 9338
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8414 994 8442
rect 966 8078 994 8106
rect 6062 8694 6090 8722
rect 2142 8302 2170 8330
rect 4998 8302 5026 8330
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 2142 8049 2170 8050
rect 2142 8023 2143 8049
rect 2143 8023 2169 8049
rect 2169 8023 2170 8049
rect 2142 8022 2170 8023
rect 6006 8022 6034 8050
rect 6566 9646 6594 9674
rect 6846 10065 6874 10066
rect 6846 10039 6847 10065
rect 6847 10039 6873 10065
rect 6873 10039 6874 10065
rect 6846 10038 6874 10039
rect 7406 10262 7434 10290
rect 6846 9897 6874 9898
rect 6846 9871 6847 9897
rect 6847 9871 6873 9897
rect 6873 9871 6874 9897
rect 6846 9870 6874 9871
rect 6510 9337 6538 9338
rect 6510 9311 6511 9337
rect 6511 9311 6537 9337
rect 6537 9311 6538 9337
rect 6510 9310 6538 9311
rect 6398 9198 6426 9226
rect 6734 9198 6762 9226
rect 6678 8918 6706 8946
rect 6902 9086 6930 9114
rect 7014 8945 7042 8946
rect 7014 8919 7015 8945
rect 7015 8919 7041 8945
rect 7041 8919 7042 8945
rect 7014 8918 7042 8919
rect 6790 8721 6818 8722
rect 6790 8695 6791 8721
rect 6791 8695 6817 8721
rect 6817 8695 6818 8721
rect 6790 8694 6818 8695
rect 7126 9198 7154 9226
rect 6566 8302 6594 8330
rect 6846 8302 6874 8330
rect 6398 8049 6426 8050
rect 6398 8023 6399 8049
rect 6399 8023 6425 8049
rect 6425 8023 6426 8049
rect 6398 8022 6426 8023
rect 2086 7966 2114 7994
rect 1022 7742 1050 7770
rect 7406 8918 7434 8946
rect 7630 9982 7658 10010
rect 8414 9870 8442 9898
rect 7630 9198 7658 9226
rect 7294 8470 7322 8498
rect 7686 8470 7714 8498
rect 7742 8385 7770 8386
rect 7742 8359 7743 8385
rect 7743 8359 7769 8385
rect 7769 8359 7770 8385
rect 7742 8358 7770 8359
rect 7126 8329 7154 8330
rect 7126 8303 7127 8329
rect 7127 8303 7153 8329
rect 7153 8303 7154 8329
rect 7126 8302 7154 8303
rect 7238 8105 7266 8106
rect 7238 8079 7239 8105
rect 7239 8079 7265 8105
rect 7265 8079 7266 8105
rect 7238 8078 7266 8079
rect 6734 7993 6762 7994
rect 6734 7967 6735 7993
rect 6735 7967 6761 7993
rect 6761 7967 6762 7993
rect 6734 7966 6762 7967
rect 7462 8022 7490 8050
rect 8806 9926 8834 9954
rect 8974 11073 9002 11074
rect 8974 11047 8975 11073
rect 8975 11047 9001 11073
rect 9001 11047 9002 11073
rect 8974 11046 9002 11047
rect 8974 10849 9002 10850
rect 8974 10823 8975 10849
rect 8975 10823 9001 10849
rect 9001 10823 9002 10849
rect 8974 10822 9002 10823
rect 8974 9897 9002 9898
rect 8974 9871 8975 9897
rect 8975 9871 9001 9897
rect 9001 9871 9002 9897
rect 8974 9870 9002 9871
rect 9646 13481 9674 13482
rect 9646 13455 9647 13481
rect 9647 13455 9673 13481
rect 9673 13455 9674 13481
rect 9646 13454 9674 13455
rect 9814 13537 9842 13538
rect 9814 13511 9815 13537
rect 9815 13511 9841 13537
rect 9841 13511 9842 13537
rect 9814 13510 9842 13511
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 10710 13174 10738 13202
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 13118 18718 13146 18746
rect 13734 18745 13762 18746
rect 13734 18719 13735 18745
rect 13735 18719 13761 18745
rect 13761 18719 13762 18745
rect 13734 18718 13762 18719
rect 11662 14041 11690 14042
rect 11662 14015 11663 14041
rect 11663 14015 11689 14041
rect 11689 14015 11690 14041
rect 11662 14014 11690 14015
rect 12110 14014 12138 14042
rect 11158 13286 11186 13314
rect 10822 13118 10850 13146
rect 9870 13089 9898 13090
rect 9870 13063 9871 13089
rect 9871 13063 9897 13089
rect 9897 13063 9898 13089
rect 9870 13062 9898 13063
rect 10654 12697 10682 12698
rect 10654 12671 10655 12697
rect 10655 12671 10681 12697
rect 10681 12671 10682 12697
rect 10654 12670 10682 12671
rect 10878 13062 10906 13090
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9254 11577 9282 11578
rect 9254 11551 9255 11577
rect 9255 11551 9281 11577
rect 9281 11551 9282 11577
rect 9254 11550 9282 11551
rect 9198 11465 9226 11466
rect 9198 11439 9199 11465
rect 9199 11439 9225 11465
rect 9225 11439 9226 11465
rect 9198 11438 9226 11439
rect 9366 11438 9394 11466
rect 9198 11158 9226 11186
rect 9198 11046 9226 11074
rect 9310 11214 9338 11242
rect 9590 11718 9618 11746
rect 9534 10990 9562 11018
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9702 11662 9730 11690
rect 9310 10934 9338 10962
rect 9086 10065 9114 10066
rect 9086 10039 9087 10065
rect 9087 10039 9113 10065
rect 9113 10039 9114 10065
rect 9086 10038 9114 10039
rect 9254 10038 9282 10066
rect 9422 10822 9450 10850
rect 9534 10793 9562 10794
rect 9534 10767 9535 10793
rect 9535 10767 9561 10793
rect 9561 10767 9562 10793
rect 9534 10766 9562 10767
rect 9926 11577 9954 11578
rect 9926 11551 9927 11577
rect 9927 11551 9953 11577
rect 9953 11551 9954 11577
rect 9926 11550 9954 11551
rect 10318 11577 10346 11578
rect 10318 11551 10319 11577
rect 10319 11551 10345 11577
rect 10345 11551 10346 11577
rect 10318 11550 10346 11551
rect 9870 11465 9898 11466
rect 9870 11439 9871 11465
rect 9871 11439 9897 11465
rect 9897 11439 9898 11465
rect 9870 11438 9898 11439
rect 9758 11158 9786 11186
rect 9870 11129 9898 11130
rect 9870 11103 9871 11129
rect 9871 11103 9897 11129
rect 9897 11103 9898 11129
rect 9870 11102 9898 11103
rect 10094 11046 10122 11074
rect 9758 10934 9786 10962
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9758 10793 9786 10794
rect 9758 10767 9759 10793
rect 9759 10767 9785 10793
rect 9785 10767 9786 10793
rect 9758 10766 9786 10767
rect 10038 10766 10066 10794
rect 9590 10038 9618 10066
rect 9142 9953 9170 9954
rect 9142 9927 9143 9953
rect 9143 9927 9169 9953
rect 9169 9927 9170 9953
rect 9142 9926 9170 9927
rect 9478 9926 9506 9954
rect 9030 9814 9058 9842
rect 9198 9870 9226 9898
rect 9030 9590 9058 9618
rect 8694 8889 8722 8890
rect 8694 8863 8695 8889
rect 8695 8863 8721 8889
rect 8721 8863 8722 8889
rect 8694 8862 8722 8863
rect 8750 8358 8778 8386
rect 7854 7966 7882 7994
rect 8526 7993 8554 7994
rect 8526 7967 8527 7993
rect 8527 7967 8553 7993
rect 8553 7967 8554 7993
rect 8526 7966 8554 7967
rect 7462 7657 7490 7658
rect 7462 7631 7463 7657
rect 7463 7631 7489 7657
rect 7489 7631 7490 7657
rect 7462 7630 7490 7631
rect 7854 7630 7882 7658
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 9254 9225 9282 9226
rect 9254 9199 9255 9225
rect 9255 9199 9281 9225
rect 9281 9199 9282 9225
rect 9254 9198 9282 9199
rect 9702 9982 9730 10010
rect 10094 10374 10122 10402
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10262 11185 10290 11186
rect 10262 11159 10263 11185
rect 10263 11159 10289 11185
rect 10289 11159 10290 11185
rect 10262 11158 10290 11159
rect 10262 11046 10290 11074
rect 10374 11662 10402 11690
rect 10486 11633 10514 11634
rect 10486 11607 10487 11633
rect 10487 11607 10513 11633
rect 10513 11607 10514 11633
rect 10486 11606 10514 11607
rect 10374 10990 10402 11018
rect 9870 9953 9898 9954
rect 9870 9927 9871 9953
rect 9871 9927 9897 9953
rect 9897 9927 9898 9953
rect 9870 9926 9898 9927
rect 10374 10374 10402 10402
rect 10318 10009 10346 10010
rect 10318 9983 10319 10009
rect 10319 9983 10345 10009
rect 10345 9983 10346 10009
rect 10318 9982 10346 9983
rect 10710 11270 10738 11298
rect 10766 11577 10794 11578
rect 10766 11551 10767 11577
rect 10767 11551 10793 11577
rect 10793 11551 10794 11577
rect 10766 11550 10794 11551
rect 10990 12697 11018 12698
rect 10990 12671 10991 12697
rect 10991 12671 11017 12697
rect 11017 12671 11018 12697
rect 10990 12670 11018 12671
rect 11158 12558 11186 12586
rect 11270 13174 11298 13202
rect 11718 13454 11746 13482
rect 11830 13201 11858 13202
rect 11830 13175 11831 13201
rect 11831 13175 11857 13201
rect 11857 13175 11858 13201
rect 11830 13174 11858 13175
rect 11494 13145 11522 13146
rect 11494 13119 11495 13145
rect 11495 13119 11521 13145
rect 11521 13119 11522 13145
rect 11494 13118 11522 13119
rect 12334 13174 12362 13202
rect 12950 13174 12978 13202
rect 12166 13062 12194 13090
rect 12670 13089 12698 13090
rect 12670 13063 12671 13089
rect 12671 13063 12697 13089
rect 12697 13063 12698 13089
rect 12670 13062 12698 13063
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 20118 17822 20146 17850
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 20118 13118 20146 13146
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 12950 12614 12978 12642
rect 12278 12558 12306 12586
rect 12222 12473 12250 12474
rect 12222 12447 12223 12473
rect 12223 12447 12249 12473
rect 12249 12447 12250 12473
rect 12222 12446 12250 12447
rect 11158 11774 11186 11802
rect 10878 11689 10906 11690
rect 10878 11663 10879 11689
rect 10879 11663 10905 11689
rect 10905 11663 10906 11689
rect 10878 11662 10906 11663
rect 10766 11214 10794 11242
rect 10990 11270 11018 11298
rect 10710 11073 10738 11074
rect 10710 11047 10711 11073
rect 10711 11047 10737 11073
rect 10737 11047 10738 11073
rect 10710 11046 10738 11047
rect 10878 10934 10906 10962
rect 10934 10401 10962 10402
rect 10934 10375 10935 10401
rect 10935 10375 10961 10401
rect 10961 10375 10962 10401
rect 10934 10374 10962 10375
rect 10710 10289 10738 10290
rect 10710 10263 10711 10289
rect 10711 10263 10737 10289
rect 10737 10263 10738 10289
rect 10710 10262 10738 10263
rect 11606 11550 11634 11578
rect 11046 11158 11074 11186
rect 11102 11073 11130 11074
rect 11102 11047 11103 11073
rect 11103 11047 11129 11073
rect 11129 11047 11130 11073
rect 11102 11046 11130 11047
rect 11214 10822 11242 10850
rect 11382 10401 11410 10402
rect 11382 10375 11383 10401
rect 11383 10375 11409 10401
rect 11409 10375 11410 10401
rect 11382 10374 11410 10375
rect 11158 10345 11186 10346
rect 11158 10319 11159 10345
rect 11159 10319 11185 10345
rect 11185 10319 11186 10345
rect 11158 10318 11186 10319
rect 10598 9926 10626 9954
rect 10038 9617 10066 9618
rect 10038 9591 10039 9617
rect 10039 9591 10065 9617
rect 10065 9591 10066 9617
rect 10038 9590 10066 9591
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9814 9337 9842 9338
rect 9814 9311 9815 9337
rect 9815 9311 9841 9337
rect 9841 9311 9842 9337
rect 9814 9310 9842 9311
rect 10150 9310 10178 9338
rect 10038 9225 10066 9226
rect 10038 9199 10039 9225
rect 10039 9199 10065 9225
rect 10065 9199 10066 9225
rect 10038 9198 10066 9199
rect 9534 9113 9562 9114
rect 9534 9087 9535 9113
rect 9535 9087 9561 9113
rect 9561 9087 9562 9113
rect 9534 9086 9562 9087
rect 9982 9113 10010 9114
rect 9982 9087 9983 9113
rect 9983 9087 10009 9113
rect 10009 9087 10010 9113
rect 9982 9086 10010 9087
rect 10318 9142 10346 9170
rect 9590 8777 9618 8778
rect 9590 8751 9591 8777
rect 9591 8751 9617 8777
rect 9617 8751 9618 8777
rect 9590 8750 9618 8751
rect 9534 8721 9562 8722
rect 9534 8695 9535 8721
rect 9535 8695 9561 8721
rect 9561 8695 9562 8721
rect 9534 8694 9562 8695
rect 10038 8694 10066 8722
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9366 8526 9394 8554
rect 9086 8497 9114 8498
rect 9086 8471 9087 8497
rect 9087 8471 9113 8497
rect 9113 8471 9114 8497
rect 9086 8470 9114 8471
rect 9030 8358 9058 8386
rect 8918 7713 8946 7714
rect 8918 7687 8919 7713
rect 8919 7687 8945 7713
rect 8945 7687 8946 7713
rect 8918 7686 8946 7687
rect 9086 8022 9114 8050
rect 10374 8862 10402 8890
rect 10430 9030 10458 9058
rect 10150 8750 10178 8778
rect 10934 9702 10962 9730
rect 10262 8470 10290 8498
rect 10542 8414 10570 8442
rect 10150 8049 10178 8050
rect 10150 8023 10151 8049
rect 10151 8023 10177 8049
rect 10177 8023 10178 8049
rect 10150 8022 10178 8023
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 8862 7294 8890 7322
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 9254 7321 9282 7322
rect 9254 7295 9255 7321
rect 9255 7295 9281 7321
rect 9281 7295 9282 7321
rect 9254 7294 9282 7295
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 11102 10121 11130 10122
rect 11102 10095 11103 10121
rect 11103 10095 11129 10121
rect 11129 10095 11130 10121
rect 11102 10094 11130 10095
rect 11438 10094 11466 10122
rect 11158 10065 11186 10066
rect 11158 10039 11159 10065
rect 11159 10039 11185 10065
rect 11185 10039 11186 10065
rect 11158 10038 11186 10039
rect 11214 9729 11242 9730
rect 11214 9703 11215 9729
rect 11215 9703 11241 9729
rect 11241 9703 11242 9729
rect 11214 9702 11242 9703
rect 10990 9198 11018 9226
rect 11102 9590 11130 9618
rect 11718 11774 11746 11802
rect 11886 11606 11914 11634
rect 11942 11550 11970 11578
rect 11718 10766 11746 10794
rect 11886 10934 11914 10962
rect 11662 10038 11690 10066
rect 11718 10318 11746 10346
rect 11270 9310 11298 9338
rect 11550 9281 11578 9282
rect 11550 9255 11551 9281
rect 11551 9255 11577 9281
rect 11577 9255 11578 9281
rect 11550 9254 11578 9255
rect 11046 8918 11074 8946
rect 10878 8833 10906 8834
rect 10878 8807 10879 8833
rect 10879 8807 10905 8833
rect 10905 8807 10906 8833
rect 10878 8806 10906 8807
rect 11438 8945 11466 8946
rect 11438 8919 11439 8945
rect 11439 8919 11465 8945
rect 11465 8919 11466 8945
rect 11438 8918 11466 8919
rect 11382 8806 11410 8834
rect 11550 8833 11578 8834
rect 11550 8807 11551 8833
rect 11551 8807 11577 8833
rect 11577 8807 11578 8833
rect 11550 8806 11578 8807
rect 10878 8441 10906 8442
rect 10878 8415 10879 8441
rect 10879 8415 10905 8441
rect 10905 8415 10906 8441
rect 10878 8414 10906 8415
rect 10766 8022 10794 8050
rect 12110 11550 12138 11578
rect 13342 12446 13370 12474
rect 13398 12614 13426 12642
rect 12614 11662 12642 11690
rect 11998 11185 12026 11186
rect 11998 11159 11999 11185
rect 11999 11159 12025 11185
rect 12025 11159 12026 11185
rect 11998 11158 12026 11159
rect 12166 11102 12194 11130
rect 11998 10318 12026 10346
rect 11718 9310 11746 9338
rect 11942 9729 11970 9730
rect 11942 9703 11943 9729
rect 11943 9703 11969 9729
rect 11969 9703 11970 9729
rect 11942 9702 11970 9703
rect 11886 9254 11914 9282
rect 11830 9086 11858 9114
rect 11718 8918 11746 8946
rect 11886 9169 11914 9170
rect 11886 9143 11887 9169
rect 11887 9143 11913 9169
rect 11913 9143 11914 9169
rect 11886 9142 11914 9143
rect 12726 11886 12754 11914
rect 12670 11633 12698 11634
rect 12670 11607 12671 11633
rect 12671 11607 12697 11633
rect 12697 11607 12698 11633
rect 12670 11606 12698 11607
rect 12950 11633 12978 11634
rect 12950 11607 12951 11633
rect 12951 11607 12977 11633
rect 12977 11607 12978 11633
rect 12950 11606 12978 11607
rect 12782 11577 12810 11578
rect 12782 11551 12783 11577
rect 12783 11551 12809 11577
rect 12809 11551 12810 11577
rect 12782 11550 12810 11551
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 13566 11913 13594 11914
rect 13566 11887 13567 11913
rect 13567 11887 13593 11913
rect 13593 11887 13594 11913
rect 13566 11886 13594 11887
rect 13230 11550 13258 11578
rect 12614 11158 12642 11186
rect 12726 11046 12754 11074
rect 12278 10934 12306 10962
rect 12166 10822 12194 10850
rect 12166 10374 12194 10402
rect 12670 10934 12698 10962
rect 12614 10793 12642 10794
rect 12614 10767 12615 10793
rect 12615 10767 12641 10793
rect 12641 10767 12642 10793
rect 12614 10766 12642 10767
rect 12894 10990 12922 11018
rect 12502 10345 12530 10346
rect 12502 10319 12503 10345
rect 12503 10319 12529 10345
rect 12529 10319 12530 10345
rect 12502 10318 12530 10319
rect 12838 10401 12866 10402
rect 12838 10375 12839 10401
rect 12839 10375 12865 10401
rect 12865 10375 12866 10401
rect 12838 10374 12866 10375
rect 12726 10318 12754 10346
rect 13118 11465 13146 11466
rect 13118 11439 13119 11465
rect 13119 11439 13145 11465
rect 13145 11439 13146 11465
rect 13118 11438 13146 11439
rect 13398 11550 13426 11578
rect 13454 11606 13482 11634
rect 13174 11102 13202 11130
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 14966 11521 14994 11522
rect 14966 11495 14967 11521
rect 14967 11495 14993 11521
rect 14993 11495 14994 11521
rect 14966 11494 14994 11495
rect 14742 11438 14770 11466
rect 13062 10934 13090 10962
rect 13286 10542 13314 10570
rect 13006 10345 13034 10346
rect 13006 10319 13007 10345
rect 13007 10319 13033 10345
rect 13033 10319 13034 10345
rect 13006 10318 13034 10319
rect 14294 11129 14322 11130
rect 14294 11103 14295 11129
rect 14295 11103 14321 11129
rect 14321 11103 14322 11129
rect 14294 11102 14322 11103
rect 14798 11102 14826 11130
rect 13622 10934 13650 10962
rect 14686 10990 14714 11018
rect 13734 10542 13762 10570
rect 13566 10374 13594 10402
rect 13454 10318 13482 10346
rect 13230 10262 13258 10290
rect 12054 9030 12082 9058
rect 11886 8806 11914 8834
rect 11886 8721 11914 8722
rect 11886 8695 11887 8721
rect 11887 8695 11913 8721
rect 11913 8695 11914 8721
rect 11886 8694 11914 8695
rect 11830 8470 11858 8498
rect 11662 8049 11690 8050
rect 11662 8023 11663 8049
rect 11663 8023 11689 8049
rect 11689 8023 11690 8049
rect 11662 8022 11690 8023
rect 13678 10289 13706 10290
rect 13678 10263 13679 10289
rect 13679 10263 13705 10289
rect 13705 10263 13706 10289
rect 13678 10262 13706 10263
rect 14294 10374 14322 10402
rect 13006 9702 13034 9730
rect 12894 9198 12922 9226
rect 14574 9617 14602 9618
rect 14574 9591 14575 9617
rect 14575 9591 14601 9617
rect 14601 9591 14602 9617
rect 14574 9590 14602 9591
rect 20006 11774 20034 11802
rect 18942 11438 18970 11466
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 20006 11102 20034 11130
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 18830 10401 18858 10402
rect 18830 10375 18831 10401
rect 18831 10375 18857 10401
rect 18857 10375 18858 10401
rect 18830 10374 18858 10375
rect 20006 10094 20034 10122
rect 13286 9225 13314 9226
rect 13286 9199 13287 9225
rect 13287 9199 13313 9225
rect 13313 9199 13314 9225
rect 13286 9198 13314 9199
rect 13622 9478 13650 9506
rect 14630 9505 14658 9506
rect 14630 9479 14631 9505
rect 14631 9479 14657 9505
rect 14657 9479 14658 9505
rect 14630 9478 14658 9479
rect 13230 8806 13258 8834
rect 12670 8526 12698 8554
rect 12782 8694 12810 8722
rect 12726 8414 12754 8442
rect 11998 8049 12026 8050
rect 11998 8023 11999 8049
rect 11999 8023 12025 8049
rect 12025 8023 12026 8049
rect 11998 8022 12026 8023
rect 10766 7657 10794 7658
rect 10766 7631 10767 7657
rect 10767 7631 10793 7657
rect 10793 7631 10794 7657
rect 10766 7630 10794 7631
rect 12222 7630 12250 7658
rect 12950 8497 12978 8498
rect 12950 8471 12951 8497
rect 12951 8471 12977 8497
rect 12977 8471 12978 8497
rect 12950 8470 12978 8471
rect 14070 9254 14098 9282
rect 13958 9142 13986 9170
rect 13342 8553 13370 8554
rect 13342 8527 13343 8553
rect 13343 8527 13369 8553
rect 13369 8527 13370 8553
rect 13342 8526 13370 8527
rect 13286 8470 13314 8498
rect 13062 8329 13090 8330
rect 13062 8303 13063 8329
rect 13063 8303 13089 8329
rect 13089 8303 13090 8329
rect 13062 8302 13090 8303
rect 13734 8441 13762 8442
rect 13734 8415 13735 8441
rect 13735 8415 13761 8441
rect 13761 8415 13762 8441
rect 13734 8414 13762 8415
rect 13566 8246 13594 8274
rect 13734 8302 13762 8330
rect 13622 8105 13650 8106
rect 13622 8079 13623 8105
rect 13623 8079 13649 8105
rect 13649 8079 13650 8105
rect 13622 8078 13650 8079
rect 13846 8078 13874 8106
rect 14798 9254 14826 9282
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 14686 9169 14714 9170
rect 14686 9143 14687 9169
rect 14687 9143 14713 9169
rect 14713 9143 14714 9169
rect 14686 9142 14714 9143
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 14406 8414 14434 8442
rect 13958 8246 13986 8274
rect 13902 7686 13930 7714
rect 12726 7657 12754 7658
rect 12726 7631 12727 7657
rect 12727 7631 12753 7657
rect 12753 7631 12754 7657
rect 12726 7630 12754 7631
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 14910 8414 14938 8442
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 18830 8134 18858 8162
rect 19950 8078 19978 8106
rect 14182 7601 14210 7602
rect 14182 7575 14183 7601
rect 14183 7575 14209 7601
rect 14209 7575 14210 7601
rect 14182 7574 14210 7575
rect 20006 7742 20034 7770
rect 18830 7574 18858 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9758 1806 9786 1834
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 10934 1833 10962 1834
rect 10934 1807 10935 1833
rect 10935 1807 10961 1833
rect 10961 1807 10962 1833
rect 10934 1806 10962 1807
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 8409 19110 8414 19138
rect 8442 19110 9030 19138
rect 9058 19110 9063 19138
rect 11769 19110 11774 19138
rect 11802 19110 12782 19138
rect 12810 19110 12815 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9417 18718 9422 18746
rect 9450 18718 10038 18746
rect 10066 18718 10071 18746
rect 13113 18718 13118 18746
rect 13146 18718 13734 18746
rect 13762 18718 13767 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 20600 17850 21000 17864
rect 20113 17822 20118 17850
rect 20146 17822 21000 17850
rect 20600 17808 21000 17822
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 11657 14014 11662 14042
rect 11690 14014 12110 14042
rect 12138 14014 12143 14042
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 6953 13510 6958 13538
rect 6986 13510 8078 13538
rect 8106 13510 8111 13538
rect 9193 13510 9198 13538
rect 9226 13510 9814 13538
rect 9842 13510 10094 13538
rect 0 13482 400 13496
rect 10066 13482 10094 13510
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 8801 13454 8806 13482
rect 8834 13454 9646 13482
rect 9674 13454 9679 13482
rect 10066 13454 11718 13482
rect 11746 13454 11751 13482
rect 0 13440 400 13454
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 11158 13314 11186 13454
rect 11153 13286 11158 13314
rect 11186 13286 11191 13314
rect 10705 13174 10710 13202
rect 10738 13174 11270 13202
rect 11298 13174 11830 13202
rect 11858 13174 12334 13202
rect 12362 13174 12950 13202
rect 12978 13174 12983 13202
rect 20600 13146 21000 13160
rect 10817 13118 10822 13146
rect 10850 13118 11494 13146
rect 11522 13118 11527 13146
rect 20113 13118 20118 13146
rect 20146 13118 21000 13146
rect 20600 13104 21000 13118
rect 9865 13062 9870 13090
rect 9898 13062 10878 13090
rect 10906 13062 10911 13090
rect 12161 13062 12166 13090
rect 12194 13062 12670 13090
rect 12698 13062 12703 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 10649 12670 10654 12698
rect 10682 12670 10990 12698
rect 11018 12670 11023 12698
rect 12945 12614 12950 12642
rect 12978 12614 13398 12642
rect 13426 12614 13431 12642
rect 11153 12558 11158 12586
rect 11186 12558 12278 12586
rect 12306 12558 12311 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 7289 12446 7294 12474
rect 7322 12446 8134 12474
rect 8162 12446 8167 12474
rect 12217 12446 12222 12474
rect 12250 12446 13342 12474
rect 13370 12446 13375 12474
rect 2137 12334 2142 12362
rect 2170 12334 5670 12362
rect 5698 12334 5703 12362
rect 6729 12278 6734 12306
rect 6762 12278 7518 12306
rect 7546 12278 7551 12306
rect 961 12222 966 12250
rect 994 12222 999 12250
rect 0 12138 400 12152
rect 966 12138 994 12222
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 0 12110 994 12138
rect 0 12096 400 12110
rect 12721 11886 12726 11914
rect 12754 11886 13566 11914
rect 13594 11886 13599 11914
rect 5665 11830 5670 11858
rect 5698 11830 7126 11858
rect 7154 11830 7159 11858
rect 20600 11802 21000 11816
rect 11153 11774 11158 11802
rect 11186 11774 11718 11802
rect 11746 11774 11751 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 9585 11718 9590 11746
rect 9618 11718 9842 11746
rect 9814 11690 9842 11718
rect 8297 11662 8302 11690
rect 8330 11662 8806 11690
rect 8834 11662 9702 11690
rect 9730 11662 9735 11690
rect 9814 11662 10374 11690
rect 10402 11662 10878 11690
rect 10906 11662 10911 11690
rect 12609 11662 12614 11690
rect 12642 11662 15974 11690
rect 7233 11606 7238 11634
rect 7266 11606 10486 11634
rect 10514 11606 11886 11634
rect 11914 11606 12670 11634
rect 12698 11606 12703 11634
rect 12945 11606 12950 11634
rect 12978 11606 13454 11634
rect 13482 11606 13487 11634
rect 15946 11578 15974 11662
rect 8969 11550 8974 11578
rect 9002 11550 9254 11578
rect 9282 11550 9287 11578
rect 9921 11550 9926 11578
rect 9954 11550 10318 11578
rect 10346 11550 10351 11578
rect 10761 11550 10766 11578
rect 10794 11550 11606 11578
rect 11634 11550 11639 11578
rect 11937 11550 11942 11578
rect 11970 11550 12110 11578
rect 12138 11550 12782 11578
rect 12810 11550 13230 11578
rect 13258 11550 13263 11578
rect 13393 11550 13398 11578
rect 13426 11522 13454 11578
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 7345 11494 7350 11522
rect 7378 11494 8190 11522
rect 8218 11494 8223 11522
rect 13426 11494 14966 11522
rect 14994 11494 14999 11522
rect 20600 11466 21000 11480
rect 8521 11438 8526 11466
rect 8554 11438 9198 11466
rect 9226 11438 9231 11466
rect 9361 11438 9366 11466
rect 9394 11438 9870 11466
rect 9898 11438 9903 11466
rect 13113 11438 13118 11466
rect 13146 11438 14742 11466
rect 14770 11438 18942 11466
rect 18970 11438 18975 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 6841 11270 6846 11298
rect 6874 11270 7070 11298
rect 7098 11270 7574 11298
rect 10705 11270 10710 11298
rect 10738 11270 10990 11298
rect 11018 11270 11023 11298
rect 7546 11242 7574 11270
rect 961 11214 966 11242
rect 994 11214 999 11242
rect 7546 11214 9310 11242
rect 9338 11214 10766 11242
rect 10794 11214 10799 11242
rect 0 11130 400 11144
rect 966 11130 994 11214
rect 2137 11158 2142 11186
rect 2170 11158 5446 11186
rect 5474 11158 6958 11186
rect 6986 11158 6991 11186
rect 7625 11158 7630 11186
rect 7658 11158 8358 11186
rect 8386 11158 8862 11186
rect 8890 11158 8895 11186
rect 9193 11158 9198 11186
rect 9226 11158 9758 11186
rect 9786 11158 10262 11186
rect 10290 11158 11046 11186
rect 11074 11158 11079 11186
rect 11993 11158 11998 11186
rect 12026 11158 12614 11186
rect 12642 11158 12647 11186
rect 15946 11158 18830 11186
rect 18858 11158 18863 11186
rect 15946 11130 15974 11158
rect 20600 11130 21000 11144
rect 0 11102 994 11130
rect 8129 11102 8134 11130
rect 8162 11102 8526 11130
rect 8554 11102 8559 11130
rect 8913 11102 8918 11130
rect 8946 11102 9870 11130
rect 9898 11102 11130 11130
rect 12161 11102 12166 11130
rect 12194 11102 13174 11130
rect 13202 11102 13454 11130
rect 14289 11102 14294 11130
rect 14322 11102 14798 11130
rect 14826 11102 15974 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 0 11088 400 11102
rect 11102 11074 11130 11102
rect 8969 11046 8974 11074
rect 9002 11046 9198 11074
rect 9226 11046 10094 11074
rect 10122 11046 10127 11074
rect 10257 11046 10262 11074
rect 10290 11046 10710 11074
rect 10738 11046 10743 11074
rect 11097 11046 11102 11074
rect 11130 11046 12726 11074
rect 12754 11046 12759 11074
rect 13426 11018 13454 11102
rect 20600 11088 21000 11102
rect 7233 10990 7238 11018
rect 7266 10990 9534 11018
rect 9562 10990 9567 11018
rect 10369 10990 10374 11018
rect 10402 10990 12894 11018
rect 12922 10990 12927 11018
rect 13426 10990 14686 11018
rect 14714 10990 14719 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 9305 10934 9310 10962
rect 9338 10934 9758 10962
rect 9786 10934 9791 10962
rect 10873 10934 10878 10962
rect 10906 10934 11886 10962
rect 11914 10934 12278 10962
rect 12306 10934 12311 10962
rect 12665 10934 12670 10962
rect 12698 10934 13062 10962
rect 13090 10934 13622 10962
rect 13650 10934 13655 10962
rect 8465 10878 8470 10906
rect 8498 10878 8806 10906
rect 8834 10878 8839 10906
rect 8969 10822 8974 10850
rect 9002 10822 9422 10850
rect 9450 10822 11214 10850
rect 11242 10822 12166 10850
rect 12194 10822 12199 10850
rect 2081 10766 2086 10794
rect 2114 10766 9534 10794
rect 9562 10766 9758 10794
rect 9786 10766 9791 10794
rect 10033 10766 10038 10794
rect 10066 10766 11718 10794
rect 11746 10766 12614 10794
rect 12642 10766 12647 10794
rect 6449 10710 6454 10738
rect 6482 10710 6902 10738
rect 6930 10710 6935 10738
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 13281 10542 13286 10570
rect 13314 10542 13734 10570
rect 13762 10542 13767 10570
rect 4186 10430 4998 10458
rect 5026 10430 6566 10458
rect 6594 10430 6599 10458
rect 4186 10402 4214 10430
rect 2137 10374 2142 10402
rect 2170 10374 4214 10402
rect 10089 10374 10094 10402
rect 10122 10374 10374 10402
rect 10402 10374 10934 10402
rect 10962 10374 10967 10402
rect 11363 10374 11382 10402
rect 11410 10374 11415 10402
rect 12161 10374 12166 10402
rect 12194 10374 12838 10402
rect 12866 10374 12871 10402
rect 13561 10374 13566 10402
rect 13594 10374 14294 10402
rect 14322 10374 18830 10402
rect 18858 10374 18863 10402
rect 11153 10318 11158 10346
rect 11186 10318 11718 10346
rect 11746 10318 11998 10346
rect 12026 10318 12502 10346
rect 12530 10318 12535 10346
rect 12721 10318 12726 10346
rect 12754 10318 13006 10346
rect 13034 10318 13454 10346
rect 13482 10318 13487 10346
rect 7401 10262 7406 10290
rect 7434 10262 10710 10290
rect 10738 10262 10743 10290
rect 13225 10262 13230 10290
rect 13258 10262 13678 10290
rect 13706 10262 13711 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 0 10122 400 10136
rect 20600 10122 21000 10136
rect 0 10094 966 10122
rect 994 10094 999 10122
rect 11097 10094 11102 10122
rect 11130 10094 11438 10122
rect 11466 10094 11471 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 0 10080 400 10094
rect 20600 10080 21000 10094
rect 6673 10038 6678 10066
rect 6706 10038 6846 10066
rect 6874 10038 6879 10066
rect 9081 10038 9086 10066
rect 9114 10038 9254 10066
rect 9282 10038 9590 10066
rect 9618 10038 9623 10066
rect 11153 10038 11158 10066
rect 11186 10038 11662 10066
rect 11690 10038 11695 10066
rect 11158 10010 11186 10038
rect 2137 9982 2142 10010
rect 2170 9982 7630 10010
rect 7658 9982 7663 10010
rect 9697 9982 9702 10010
rect 9730 9982 10318 10010
rect 10346 9982 11186 10010
rect 8801 9926 8806 9954
rect 8834 9926 9142 9954
rect 9170 9926 9175 9954
rect 9473 9926 9478 9954
rect 9506 9926 9870 9954
rect 9898 9926 10598 9954
rect 10626 9926 10631 9954
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 6057 9870 6062 9898
rect 6090 9870 6846 9898
rect 6874 9870 6879 9898
rect 8409 9870 8414 9898
rect 8442 9870 8974 9898
rect 9002 9870 9198 9898
rect 9226 9870 9231 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 9025 9814 9030 9842
rect 9058 9814 9063 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 0 9758 994 9786
rect 0 9744 400 9758
rect 4186 9646 4998 9674
rect 5026 9646 6566 9674
rect 6594 9646 6599 9674
rect 4186 9618 4214 9646
rect 9030 9618 9058 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 10929 9702 10934 9730
rect 10962 9702 11214 9730
rect 11242 9702 11382 9730
rect 11410 9702 11415 9730
rect 11937 9702 11942 9730
rect 11970 9702 13006 9730
rect 13034 9702 13454 9730
rect 13426 9618 13454 9702
rect 2137 9590 2142 9618
rect 2170 9590 4214 9618
rect 9025 9590 9030 9618
rect 9058 9590 9063 9618
rect 10033 9590 10038 9618
rect 10066 9590 11102 9618
rect 11130 9590 11135 9618
rect 13426 9590 14574 9618
rect 14602 9590 14607 9618
rect 13617 9478 13622 9506
rect 13650 9478 14630 9506
rect 14658 9478 14663 9506
rect 0 9450 400 9464
rect 0 9422 966 9450
rect 994 9422 999 9450
rect 0 9408 400 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 5833 9310 5838 9338
rect 5866 9310 6510 9338
rect 6538 9310 6543 9338
rect 9809 9310 9814 9338
rect 9842 9310 10150 9338
rect 10178 9310 10183 9338
rect 11265 9310 11270 9338
rect 11298 9310 11718 9338
rect 11746 9310 11751 9338
rect 11545 9254 11550 9282
rect 11578 9254 11886 9282
rect 11914 9254 11919 9282
rect 14065 9254 14070 9282
rect 14098 9254 14798 9282
rect 14826 9254 14831 9282
rect 6393 9198 6398 9226
rect 6426 9198 6734 9226
rect 6762 9198 7126 9226
rect 7154 9198 7159 9226
rect 7625 9198 7630 9226
rect 7658 9198 9254 9226
rect 9282 9198 9287 9226
rect 10033 9198 10038 9226
rect 10066 9198 10990 9226
rect 11018 9198 11023 9226
rect 12889 9198 12894 9226
rect 12922 9198 13286 9226
rect 13314 9198 13319 9226
rect 15946 9198 18830 9226
rect 18858 9198 18863 9226
rect 15946 9170 15974 9198
rect 10313 9142 10318 9170
rect 10346 9142 11886 9170
rect 11914 9142 11919 9170
rect 13953 9142 13958 9170
rect 13986 9142 14686 9170
rect 14714 9142 15974 9170
rect 20600 9114 21000 9128
rect 6897 9086 6902 9114
rect 6930 9086 9534 9114
rect 9562 9086 9567 9114
rect 9977 9086 9982 9114
rect 10010 9086 11830 9114
rect 11858 9086 11863 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 10425 9030 10430 9058
rect 10458 9030 12054 9058
rect 12082 9030 12087 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 6673 8918 6678 8946
rect 6706 8918 7014 8946
rect 7042 8918 7406 8946
rect 7434 8918 7439 8946
rect 11041 8918 11046 8946
rect 11074 8918 11438 8946
rect 11466 8918 11718 8946
rect 11746 8918 11751 8946
rect 8689 8862 8694 8890
rect 8722 8862 10374 8890
rect 10402 8862 10407 8890
rect 10873 8806 10878 8834
rect 10906 8806 11382 8834
rect 11410 8806 11550 8834
rect 11578 8806 11583 8834
rect 11881 8806 11886 8834
rect 11914 8806 13230 8834
rect 13258 8806 13263 8834
rect 9585 8750 9590 8778
rect 9618 8750 10150 8778
rect 10178 8750 10183 8778
rect 6057 8694 6062 8722
rect 6090 8694 6790 8722
rect 6818 8694 6823 8722
rect 9529 8694 9534 8722
rect 9562 8694 10038 8722
rect 10066 8694 10071 8722
rect 11881 8694 11886 8722
rect 11914 8694 12782 8722
rect 12810 8694 12815 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7686 8526 9366 8554
rect 9394 8526 9399 8554
rect 12665 8526 12670 8554
rect 12698 8526 13342 8554
rect 13370 8526 13375 8554
rect 7686 8498 7714 8526
rect 7289 8470 7294 8498
rect 7322 8470 7686 8498
rect 7714 8470 7719 8498
rect 9081 8470 9086 8498
rect 9114 8470 10262 8498
rect 10290 8470 10295 8498
rect 11825 8470 11830 8498
rect 11858 8470 12950 8498
rect 12978 8470 12983 8498
rect 13281 8470 13286 8498
rect 13314 8470 13319 8498
rect 0 8442 400 8456
rect 13286 8442 13314 8470
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 10537 8414 10542 8442
rect 10570 8414 10878 8442
rect 10906 8414 10911 8442
rect 12721 8414 12726 8442
rect 12754 8414 13734 8442
rect 13762 8414 14406 8442
rect 14434 8414 14910 8442
rect 14938 8414 14943 8442
rect 0 8400 400 8414
rect 7546 8358 7742 8386
rect 7770 8358 7775 8386
rect 8745 8358 8750 8386
rect 8778 8358 9030 8386
rect 9058 8358 9063 8386
rect 7546 8330 7574 8358
rect 2137 8302 2142 8330
rect 2170 8302 4998 8330
rect 5026 8302 6566 8330
rect 6594 8302 6846 8330
rect 6874 8302 6879 8330
rect 7121 8302 7126 8330
rect 7154 8302 7574 8330
rect 13057 8302 13062 8330
rect 13090 8302 13734 8330
rect 13762 8302 13767 8330
rect 13561 8246 13566 8274
rect 13594 8246 13958 8274
rect 13986 8246 13991 8274
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 15946 8134 18830 8162
rect 18858 8134 18863 8162
rect 0 8106 400 8120
rect 15946 8106 15974 8134
rect 20600 8106 21000 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 6006 8078 7238 8106
rect 7266 8078 7271 8106
rect 13617 8078 13622 8106
rect 13650 8078 13846 8106
rect 13874 8078 15974 8106
rect 19945 8078 19950 8106
rect 19978 8078 21000 8106
rect 0 8064 400 8078
rect 6006 8050 6034 8078
rect 20600 8064 21000 8078
rect 2137 8022 2142 8050
rect 2170 8022 6006 8050
rect 6034 8022 6039 8050
rect 6393 8022 6398 8050
rect 6426 8022 7462 8050
rect 7490 8022 9086 8050
rect 9114 8022 9119 8050
rect 10145 8022 10150 8050
rect 10178 8022 10766 8050
rect 10794 8022 10799 8050
rect 11657 8022 11662 8050
rect 11690 8022 11998 8050
rect 12026 8022 12031 8050
rect 10150 7994 10178 8022
rect 2081 7966 2086 7994
rect 2114 7966 6734 7994
rect 6762 7966 6767 7994
rect 7849 7966 7854 7994
rect 7882 7966 8526 7994
rect 8554 7966 10178 7994
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 0 7770 400 7784
rect 20600 7770 21000 7784
rect 0 7742 1022 7770
rect 1050 7742 1055 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 0 7728 400 7742
rect 20600 7728 21000 7742
rect 8913 7686 8918 7714
rect 8946 7686 13902 7714
rect 13930 7686 13935 7714
rect 7457 7630 7462 7658
rect 7490 7630 7854 7658
rect 7882 7630 7887 7658
rect 10761 7630 10766 7658
rect 10794 7630 12222 7658
rect 12250 7630 12726 7658
rect 12754 7630 12759 7658
rect 14177 7574 14182 7602
rect 14210 7574 18830 7602
rect 18858 7574 18863 7602
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 8857 7294 8862 7322
rect 8890 7294 9254 7322
rect 9282 7294 9287 7322
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 9753 1806 9758 1834
rect 9786 1806 10934 1834
rect 10962 1806 10967 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 11382 10374 11410 10402
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 11382 9702 11410 9730
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 11382 10402 11410 10407
rect 11382 9730 11410 10374
rect 11382 9697 11410 9702
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _091_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10024 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _092_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _093_
timestamp 1698175906
transform -1 0 11760 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _094_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11200 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _095_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 -1 10192
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6832 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8288 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1698175906
transform 1 0 8736 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform 1 0 9072 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _100_
timestamp 1698175906
transform 1 0 10248 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6776 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7000 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _103_
timestamp 1698175906
transform 1 0 8904 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1698175906
transform 1 0 8960 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9912 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform 1 0 9072 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform -1 0 11368 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _108_
timestamp 1698175906
transform 1 0 10808 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11648 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _111_
timestamp 1698175906
transform -1 0 8960 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _112_
timestamp 1698175906
transform 1 0 11312 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11480 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11480 0 -1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _115_
timestamp 1698175906
transform -1 0 11368 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _116_
timestamp 1698175906
transform -1 0 11032 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _117_
timestamp 1698175906
transform -1 0 10248 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform -1 0 10136 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _119_
timestamp 1698175906
transform -1 0 9352 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _120_
timestamp 1698175906
transform 1 0 8736 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8064 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 10136 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _123_
timestamp 1698175906
transform -1 0 9800 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform 1 0 12768 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform -1 0 12824 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 8736 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform 1 0 14000 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _128_
timestamp 1698175906
transform 1 0 13160 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698175906
transform -1 0 12096 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 10640 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _131_
timestamp 1698175906
transform -1 0 12768 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13216 0 -1 11760
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1698175906
transform 1 0 13496 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform -1 0 12096 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform 1 0 11648 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _136_
timestamp 1698175906
transform -1 0 14000 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13160 0 -1 8624
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 8736 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _139_
timestamp 1698175906
transform -1 0 8344 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 12432 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11592 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 13832 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _143_
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 9016 0 -1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _145_
timestamp 1698175906
transform 1 0 8344 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform -1 0 11816 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _147_
timestamp 1698175906
transform 1 0 10584 0 -1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform 1 0 11424 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _149_
timestamp 1698175906
transform -1 0 11312 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1698175906
transform -1 0 10472 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12320 0 1 10192
box -43 -43 1051 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _152_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11480 0 1 10976
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _153_
timestamp 1698175906
transform -1 0 11928 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _154_
timestamp 1698175906
transform -1 0 11256 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 11256 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _156_
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _157_
timestamp 1698175906
transform -1 0 14392 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _158_
timestamp 1698175906
transform -1 0 13776 0 1 10976
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _159_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11928 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _160_
timestamp 1698175906
transform -1 0 12768 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform 1 0 13440 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _162_
timestamp 1698175906
transform -1 0 13272 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _163_
timestamp 1698175906
transform 1 0 6944 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _164_
timestamp 1698175906
transform 1 0 7392 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _165_
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9800 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _167_
timestamp 1698175906
transform -1 0 7392 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _168_
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _170_
timestamp 1698175906
transform 1 0 6328 0 -1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _171_
timestamp 1698175906
transform 1 0 5768 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform 1 0 6440 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _173_
timestamp 1698175906
transform -1 0 7448 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform -1 0 7000 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _175_
timestamp 1698175906
transform 1 0 9240 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _176_
timestamp 1698175906
transform 1 0 9912 0 -1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _177_
timestamp 1698175906
transform 1 0 9352 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _178_
timestamp 1698175906
transform 1 0 9800 0 1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _179_
timestamp 1698175906
transform -1 0 7336 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _180_
timestamp 1698175906
transform 1 0 7616 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _181_
timestamp 1698175906
transform 1 0 6776 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7000 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _183_
timestamp 1698175906
transform 1 0 8008 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _184_
timestamp 1698175906
transform 1 0 10640 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _185_
timestamp 1698175906
transform 1 0 9016 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _186_
timestamp 1698175906
transform 1 0 6888 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _187_
timestamp 1698175906
transform 1 0 8904 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _188_
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _189_
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _190_
timestamp 1698175906
transform 1 0 12096 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _191_
timestamp 1698175906
transform 1 0 6832 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_
timestamp 1698175906
transform 1 0 13160 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform 1 0 7728 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 11200 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform -1 0 11424 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform 1 0 13272 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 11872 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 12768 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform -1 0 7224 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform -1 0 6552 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform -1 0 6552 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform -1 0 6552 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform -1 0 9184 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform -1 0 7616 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698175906
transform -1 0 7000 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12376 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__CLK
timestamp 1698175906
transform 1 0 14392 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__CLK
timestamp 1698175906
transform 1 0 14952 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__CLK
timestamp 1698175906
transform 1 0 13720 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 14896 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 12320 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 12936 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 11816 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 13608 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 15064 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9520 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_120 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_124 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7616 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_126 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7728 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_131
timestamp 1698175906
transform 1 0 8008 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698175906
transform 1 0 8232 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 11760 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 11984 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 12208 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 12208 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_125
timestamp 1698175906
transform 1 0 7672 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_155
timestamp 1698175906
transform 1 0 9352 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_193 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11480 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_201
timestamp 1698175906
transform 1 0 11928 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_205
timestamp 1698175906
transform 1 0 12152 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_209
timestamp 1698175906
transform 1 0 12376 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 14168 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698175906
transform 1 0 5600 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_92
timestamp 1698175906
transform 1 0 5824 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_94
timestamp 1698175906
transform 1 0 5936 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_124
timestamp 1698175906
transform 1 0 7616 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 12264 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 12376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_243
timestamp 1698175906
transform 1 0 14280 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_247
timestamp 1698175906
transform 1 0 14504 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 16296 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 2464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_69
timestamp 1698175906
transform 1 0 4536 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_73
timestamp 1698175906
transform 1 0 4760 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_75
timestamp 1698175906
transform 1 0 4872 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_113
timestamp 1698175906
transform 1 0 7000 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_119
timestamp 1698175906
transform 1 0 7336 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_135
timestamp 1698175906
transform 1 0 8232 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_145
timestamp 1698175906
transform 1 0 8792 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_161
timestamp 1698175906
transform 1 0 9688 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_165
timestamp 1698175906
transform 1 0 9912 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 10248 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 11032 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698175906
transform 1 0 11256 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_191
timestamp 1698175906
transform 1 0 11368 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 14280 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_108
timestamp 1698175906
transform 1 0 6720 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_119
timestamp 1698175906
transform 1 0 7336 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_123
timestamp 1698175906
transform 1 0 7560 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_130
timestamp 1698175906
transform 1 0 7952 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_171
timestamp 1698175906
transform 1 0 10248 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_179
timestamp 1698175906
transform 1 0 10696 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_187
timestamp 1698175906
transform 1 0 11144 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_189
timestamp 1698175906
transform 1 0 11256 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_194
timestamp 1698175906
transform 1 0 11536 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_231
timestamp 1698175906
transform 1 0 13608 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_235
timestamp 1698175906
transform 1 0 13832 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_267
timestamp 1698175906
transform 1 0 15624 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698175906
transform 1 0 16072 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_117
timestamp 1698175906
transform 1 0 7224 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_121
timestamp 1698175906
transform 1 0 7448 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_152
timestamp 1698175906
transform 1 0 9184 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_154
timestamp 1698175906
transform 1 0 9296 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_202
timestamp 1698175906
transform 1 0 11984 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_234
timestamp 1698175906
transform 1 0 13776 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_240
timestamp 1698175906
transform 1 0 14112 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_90
timestamp 1698175906
transform 1 0 5712 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_95
timestamp 1698175906
transform 1 0 5992 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_99
timestamp 1698175906
transform 1 0 6216 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_111
timestamp 1698175906
transform 1 0 6888 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_113
timestamp 1698175906
transform 1 0 7000 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_120
timestamp 1698175906
transform 1 0 7392 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 8288 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_152
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_164
timestamp 1698175906
transform 1 0 9856 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_177
timestamp 1698175906
transform 1 0 10584 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_179
timestamp 1698175906
transform 1 0 10696 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_202
timestamp 1698175906
transform 1 0 11984 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698175906
transform 1 0 12992 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_222
timestamp 1698175906
transform 1 0 13104 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_252
timestamp 1698175906
transform 1 0 14784 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_256
timestamp 1698175906
transform 1 0 15008 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_272
timestamp 1698175906
transform 1 0 15904 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 4760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 4872 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_109
timestamp 1698175906
transform 1 0 6776 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_116
timestamp 1698175906
transform 1 0 7168 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_132
timestamp 1698175906
transform 1 0 8064 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_140
timestamp 1698175906
transform 1 0 8512 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_169
timestamp 1698175906
transform 1 0 10136 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_177
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_185
timestamp 1698175906
transform 1 0 11032 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_191
timestamp 1698175906
transform 1 0 11368 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_202
timestamp 1698175906
transform 1 0 11984 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_210
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_214
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_255
timestamp 1698175906
transform 1 0 14952 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_259
timestamp 1698175906
transform 1 0 15176 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_291
timestamp 1698175906
transform 1 0 16968 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_307
timestamp 1698175906
transform 1 0 17864 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_88
timestamp 1698175906
transform 1 0 5600 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_96
timestamp 1698175906
transform 1 0 6048 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_100
timestamp 1698175906
transform 1 0 6272 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_102
timestamp 1698175906
transform 1 0 6384 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_113
timestamp 1698175906
transform 1 0 7000 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_129
timestamp 1698175906
transform 1 0 7896 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_137
timestamp 1698175906
transform 1 0 8344 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 8456 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_146
timestamp 1698175906
transform 1 0 8848 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_167
timestamp 1698175906
transform 1 0 10024 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_175
timestamp 1698175906
transform 1 0 10472 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_183
timestamp 1698175906
transform 1 0 10920 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_189
timestamp 1698175906
transform 1 0 11256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_197
timestamp 1698175906
transform 1 0 11704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_204
timestamp 1698175906
transform 1 0 12096 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698175906
transform 1 0 12320 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_254
timestamp 1698175906
transform 1 0 14896 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_258
timestamp 1698175906
transform 1 0 15120 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_113
timestamp 1698175906
transform 1 0 7000 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_121
timestamp 1698175906
transform 1 0 7448 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_222
timestamp 1698175906
transform 1 0 13104 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_226
timestamp 1698175906
transform 1 0 13328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_233
timestamp 1698175906
transform 1 0 13720 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 14168 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_121
timestamp 1698175906
transform 1 0 7448 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_129
timestamp 1698175906
transform 1 0 7896 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_133
timestamp 1698175906
transform 1 0 8120 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_135
timestamp 1698175906
transform 1 0 8232 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_156
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_262
timestamp 1698175906
transform 1 0 15344 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_117
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_125
timestamp 1698175906
transform 1 0 7672 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_129
timestamp 1698175906
transform 1 0 7896 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_131
timestamp 1698175906
transform 1 0 8008 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_140
timestamp 1698175906
transform 1 0 8512 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_184
timestamp 1698175906
transform 1 0 10976 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_191
timestamp 1698175906
transform 1 0 11368 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_210
timestamp 1698175906
transform 1 0 12432 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_218
timestamp 1698175906
transform 1 0 12880 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_234
timestamp 1698175906
transform 1 0 13776 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_238
timestamp 1698175906
transform 1 0 14000 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_240
timestamp 1698175906
transform 1 0 14112 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1698175906
transform 1 0 6496 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_108
timestamp 1698175906
transform 1 0 6720 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_110
timestamp 1698175906
transform 1 0 6832 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_155
timestamp 1698175906
transform 1 0 9352 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_167
timestamp 1698175906
transform 1 0 10024 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_190
timestamp 1698175906
transform 1 0 11312 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_194
timestamp 1698175906
transform 1 0 11536 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_201
timestamp 1698175906
transform 1 0 11928 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 12376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_253
timestamp 1698175906
transform 1 0 14840 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_257
timestamp 1698175906
transform 1 0 15064 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 15960 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_111
timestamp 1698175906
transform 1 0 6888 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_126
timestamp 1698175906
transform 1 0 7728 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_142
timestamp 1698175906
transform 1 0 8624 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_150
timestamp 1698175906
transform 1 0 9072 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_154
timestamp 1698175906
transform 1 0 9296 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698175906
transform 1 0 9800 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 10248 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698175906
transform 1 0 11032 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_187
timestamp 1698175906
transform 1 0 11144 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_217
timestamp 1698175906
transform 1 0 12824 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_221
timestamp 1698175906
transform 1 0 13048 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_233
timestamp 1698175906
transform 1 0 13720 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 4032 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_117
timestamp 1698175906
transform 1 0 7224 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_125
timestamp 1698175906
transform 1 0 7672 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_137
timestamp 1698175906
transform 1 0 8344 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_146
timestamp 1698175906
transform 1 0 8848 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_176
timestamp 1698175906
transform 1 0 10528 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_192
timestamp 1698175906
transform 1 0 11424 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_200
timestamp 1698175906
transform 1 0 11872 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 16128 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698175906
transform 1 0 6776 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_144
timestamp 1698175906
transform 1 0 8736 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_154
timestamp 1698175906
transform 1 0 9296 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_170
timestamp 1698175906
transform 1 0 10192 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_189
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698175906
transform 1 0 11704 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_199
timestamp 1698175906
transform 1 0 11816 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_229
timestamp 1698175906
transform 1 0 13496 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_233
timestamp 1698175906
transform 1 0 13720 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 14168 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 8288 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_148
timestamp 1698175906
transform 1 0 8960 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_156
timestamp 1698175906
transform 1 0 9408 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_160
timestamp 1698175906
transform 1 0 9632 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_162
timestamp 1698175906
transform 1 0 9744 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_197
timestamp 1698175906
transform 1 0 11704 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_201
timestamp 1698175906
transform 1 0 11928 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_216
timestamp 1698175906
transform 1 0 12768 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_165
timestamp 1698175906
transform 1 0 9912 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 10360 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_206
timestamp 1698175906
transform 1 0 12208 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_210
timestamp 1698175906
transform 1 0 12432 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_333
timestamp 1698175906
transform 1 0 19320 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_341
timestamp 1698175906
transform 1 0 19768 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_174
timestamp 1698175906
transform 1 0 10416 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_190
timestamp 1698175906
transform 1 0 11312 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_199
timestamp 1698175906
transform 1 0 11816 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 12264 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698175906
transform 1 0 19320 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_341
timestamp 1698175906
transform 1 0 19768 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_156
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_183
timestamp 1698175906
transform 1 0 10920 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_199
timestamp 1698175906
transform 1 0 11816 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_220
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_222
timestamp 1698175906
transform 1 0 13104 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_249
timestamp 1698175906
transform 1 0 14616 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_265
timestamp 1698175906
transform 1 0 15512 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_273
timestamp 1698175906
transform 1 0 15960 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1698175906
transform 1 0 16184 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_169
timestamp 1698175906
transform 1 0 10136 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita36_23 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10136 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita36_24
timestamp 1698175906
transform 1 0 19992 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita36_25
timestamp 1698175906
transform -1 0 8008 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita36_26
timestamp 1698175906
transform 1 0 19992 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 2240 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 2240 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 2240 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 8456 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 9464 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform -1 0 2240 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 13160 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 7728 400 7784 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 17808 21000 17864 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 7728 0 7784 400 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 9408 400 9464 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 10080 400 10136 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 11760 20600 11816 21000 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 12096 400 12152 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 11088 400 11144 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 13104 20600 13160 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 7532 12152 7532 12152 0 _000_
rlabel metal2 6076 8400 6076 8400 0 _001_
rlabel metal2 5908 9436 5908 9436 0 _002_
rlabel metal3 6468 9884 6468 9884 0 _003_
rlabel metal3 9548 8876 9548 8876 0 _004_
rlabel metal3 9688 8484 9688 8484 0 _005_
rlabel metal2 7140 7868 7140 7868 0 _006_
rlabel metal2 6748 10612 6748 10612 0 _007_
rlabel metal2 8484 13454 8484 13454 0 _008_
rlabel metal2 11452 8008 11452 8008 0 _009_
rlabel metal2 9492 7812 9492 7812 0 _010_
rlabel metal2 8204 11368 8204 11368 0 _011_
rlabel metal2 9660 12152 9660 12152 0 _012_
rlabel metal2 13216 7700 13216 7700 0 _013_
rlabel metal2 13664 11620 13664 11620 0 _014_
rlabel metal2 12572 8316 12572 8316 0 _015_
rlabel metal2 7308 12572 7308 12572 0 _016_
rlabel metal2 13636 9352 13636 9352 0 _017_
rlabel metal2 8204 7434 8204 7434 0 _018_
rlabel metal2 11256 13468 11256 13468 0 _019_
rlabel metal2 11676 11704 11676 11704 0 _020_
rlabel metal2 10948 12964 10948 12964 0 _021_
rlabel metal2 13748 10304 13748 10304 0 _022_
rlabel metal2 12348 12908 12348 12908 0 _023_
rlabel metal2 13244 9688 13244 9688 0 _024_
rlabel metal2 14700 10304 14700 10304 0 _025_
rlabel metal3 14014 9604 14014 9604 0 _026_
rlabel metal2 14084 9044 14084 9044 0 _027_
rlabel metal2 8764 7896 8764 7896 0 _028_
rlabel metal2 11564 13580 11564 13580 0 _029_
rlabel metal2 10864 12684 10864 12684 0 _030_
rlabel metal2 11732 12012 11732 12012 0 _031_
rlabel metal3 11424 10052 11424 10052 0 _032_
rlabel metal2 11760 11172 11760 11172 0 _033_
rlabel metal2 11844 11256 11844 11256 0 _034_
rlabel metal2 10752 12628 10752 12628 0 _035_
rlabel metal3 10836 12684 10836 12684 0 _036_
rlabel metal2 13972 11172 13972 11172 0 _037_
rlabel metal2 12180 12768 12180 12768 0 _038_
rlabel metal2 13244 10136 13244 10136 0 _039_
rlabel metal2 7280 11956 7280 11956 0 _040_
rlabel metal2 6636 8568 6636 8568 0 _041_
rlabel metal2 7308 8848 7308 8848 0 _042_
rlabel metal2 6412 9380 6412 9380 0 _043_
rlabel metal2 7420 10528 7420 10528 0 _044_
rlabel metal2 5852 9268 5852 9268 0 _045_
rlabel metal3 6776 10052 6776 10052 0 _046_
rlabel metal2 7308 10402 7308 10402 0 _047_
rlabel metal2 10164 9296 10164 9296 0 _048_
rlabel metal2 10052 8736 10052 8736 0 _049_
rlabel metal2 7196 8176 7196 8176 0 _050_
rlabel metal3 7350 8316 7350 8316 0 _051_
rlabel metal2 9240 10780 9240 10780 0 _052_
rlabel metal2 9436 10416 9436 10416 0 _053_
rlabel metal2 10892 9044 10892 9044 0 _054_
rlabel metal3 10248 9940 10248 9940 0 _055_
rlabel metal2 6916 9380 6916 9380 0 _056_
rlabel metal2 6804 10360 6804 10360 0 _057_
rlabel metal3 9100 9884 9100 9884 0 _058_
rlabel metal2 10388 10220 10388 10220 0 _059_
rlabel metal2 6860 11228 6860 11228 0 _060_
rlabel metal2 7252 11732 7252 11732 0 _061_
rlabel metal2 6888 10500 6888 10500 0 _062_
rlabel metal2 8848 12684 8848 12684 0 _063_
rlabel metal2 11732 13692 11732 13692 0 _064_
rlabel metal3 9240 13468 9240 13468 0 _065_
rlabel metal3 10668 11172 10668 11172 0 _066_
rlabel metal3 11928 11060 11928 11060 0 _067_
rlabel metal2 11340 9380 11340 9380 0 _068_
rlabel metal2 10052 9856 10052 9856 0 _069_
rlabel metal2 7252 10892 7252 10892 0 _070_
rlabel metal2 12012 10192 12012 10192 0 _071_
rlabel metal2 11900 8988 11900 8988 0 _072_
rlabel metal3 11312 9716 11312 9716 0 _073_
rlabel metal3 10472 8036 10472 8036 0 _074_
rlabel metal2 9828 9492 9828 9492 0 _075_
rlabel metal3 8344 11116 8344 11116 0 _076_
rlabel metal2 7644 12152 7644 12152 0 _077_
rlabel metal3 10360 11676 10360 11676 0 _078_
rlabel metal2 13468 11368 13468 11368 0 _079_
rlabel metal2 12684 9156 12684 9156 0 _080_
rlabel metal2 13916 7840 13916 7840 0 _081_
rlabel metal2 14140 8204 14140 8204 0 _082_
rlabel metal3 12376 11564 12376 11564 0 _083_
rlabel metal2 10892 10724 10892 10724 0 _084_
rlabel metal2 13636 11060 13636 11060 0 _085_
rlabel metal2 12740 11788 12740 11788 0 _086_
rlabel metal2 11844 8232 11844 8232 0 _087_
rlabel metal3 12348 8708 12348 8708 0 _088_
rlabel metal2 13748 8176 13748 8176 0 _089_
rlabel metal2 8316 12488 8316 12488 0 _090_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 11732 10752 11732 10752 0 clknet_0_clk
rlabel metal2 6972 13132 6972 13132 0 clknet_1_0__leaf_clk
rlabel metal2 15008 11508 15008 11508 0 clknet_1_1__leaf_clk
rlabel metal3 11844 8036 11844 8036 0 dut36.count\[0\]
rlabel metal3 10724 8428 10724 8428 0 dut36.count\[1\]
rlabel metal2 8372 10864 8372 10864 0 dut36.count\[2\]
rlabel metal3 10500 11060 10500 11060 0 dut36.count\[3\]
rlabel metal2 14812 10528 14812 10528 0 net1
rlabel metal3 3178 10388 3178 10388 0 net10
rlabel metal3 11900 14028 11900 14028 0 net11
rlabel metal2 13580 10360 13580 10360 0 net12
rlabel metal2 5684 12320 5684 12320 0 net13
rlabel metal2 8820 2982 8820 2982 0 net14
rlabel metal2 13972 8960 13972 8960 0 net15
rlabel metal2 8484 15960 8484 15960 0 net16
rlabel metal2 13860 8036 13860 8036 0 net17
rlabel metal2 14756 11480 14756 11480 0 net18
rlabel metal2 14168 7924 14168 7924 0 net19
rlabel metal2 7644 9436 7644 9436 0 net2
rlabel metal2 9772 13524 9772 13524 0 net20
rlabel metal2 5460 10948 5460 10948 0 net21
rlabel metal2 13384 12796 13384 12796 0 net22
rlabel metal2 9996 19376 9996 19376 0 net23
rlabel metal2 20132 17976 20132 17976 0 net24
rlabel metal2 7756 1015 7756 1015 0 net25
rlabel metal2 20132 13272 20132 13272 0 net26
rlabel metal2 10388 2982 10388 2982 0 net3
rlabel metal2 6048 7588 6048 7588 0 net4
rlabel metal2 2100 8204 2100 8204 0 net5
rlabel metal2 2156 8568 2156 8568 0 net6
rlabel metal3 15960 11620 15960 11620 0 net7
rlabel metal2 10976 13188 10976 13188 0 net8
rlabel metal3 3178 9604 3178 9604 0 net9
rlabel metal2 20020 11172 20020 11172 0 segm[10]
rlabel metal3 679 9772 679 9772 0 segm[11]
rlabel metal2 9772 1099 9772 1099 0 segm[12]
rlabel metal3 707 7756 707 7756 0 segm[13]
rlabel metal3 679 8092 679 8092 0 segm[1]
rlabel metal3 679 8428 679 8428 0 segm[4]
rlabel metal3 20321 11452 20321 11452 0 segm[6]
rlabel metal2 11116 19873 11116 19873 0 segm[7]
rlabel metal3 679 9436 679 9436 0 segm[8]
rlabel metal3 679 10108 679 10108 0 segm[9]
rlabel metal2 11788 19873 11788 19873 0 sel[0]
rlabel metal2 20020 10276 20020 10276 0 sel[10]
rlabel metal3 679 12124 679 12124 0 sel[11]
rlabel metal2 9100 1099 9100 1099 0 sel[1]
rlabel metal3 20321 9100 20321 9100 0 sel[2]
rlabel metal2 8428 19873 8428 19873 0 sel[3]
rlabel metal2 19964 8232 19964 8232 0 sel[4]
rlabel metal2 20020 11900 20020 11900 0 sel[5]
rlabel metal2 20020 7924 20020 7924 0 sel[6]
rlabel metal3 9744 18732 9744 18732 0 sel[7]
rlabel metal3 679 11116 679 11116 0 sel[8]
rlabel metal2 13132 19677 13132 19677 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
